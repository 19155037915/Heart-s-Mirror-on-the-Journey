`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/10/23 22:25:17
// Design Name: 
// Module Name: ui_display
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


// ui_display.v

module ui_display(
    input             lcd_pclk,      // lcd驱动时钟
    input             sys_rst_n,     // 复位信号
    
    input      [31:0] touch_data,    // 触摸坐标数据
    input      [1:0]  ui_state,      // 界面状态
    input      [2:0]   data_state,
    input      [2:0]   data_sel  ,

    //ADC数据显示
    input      [15:0] xinlv_bcd,
    input      [15:0] hrv_bcd,
    input      [1:0] arrhythmia_level,
    input      [15:0] rr_bcd,
    
    input      [10:0] pixel_xpos,    // 像素点横坐标
    input      [10:0] pixel_ypos,    // 像素点纵坐标
    output reg [23:0] pixel_data     // 像素点数据
);

//wire define
wire   [3:0]              xinlv_bcd_1    ;  // 心率个位数
wire   [3:0]              xinlv_bcd_2    ;  // 心率十位数
wire   [3:0]              xinlv_bcd_3    ;  // 心率百位数

wire   [3:0]              rr_bcd_1    ;  // RR个位数
wire   [3:0]              rr_bcd_2    ;  // RR十位数
wire   [3:0]              rr_bcd_3    ;  // RR百位数

wire   [3:0]              hrv_bcd_1    ;  // hrv个位数
wire   [3:0]              hrv_bcd_2    ;  // hrv十位数
wire   [3:0]              hrv_bcd_3    ;  // hrv百位数

//赋值
assign  xinlv_bcd_1 = xinlv_bcd[11:8] ;   // 心率百位数
assign  xinlv_bcd_2 = xinlv_bcd[7:4] ;   // 心率十位数
assign  xinlv_bcd_3 = xinlv_bcd[3:0] ;   // 心率个位数

assign  rr_bcd_1 = rr_bcd[11:8] ;   // RR百位数
assign  rr_bcd_2 = rr_bcd[7:4] ;   // RR十位数
assign  rr_bcd_3 = rr_bcd[3:0] ;   // RR个位数

assign  hrv_bcd_1 = hrv_bcd[11:8] ;   // hrv百位数
assign  hrv_bcd_2 = hrv_bcd[7:4] ;   // hrv十位数
assign  hrv_bcd_3 = hrv_bcd[3:0] ;   // hrv个位数

//状态显示
reg [5:0] level_state [3:0];

always@(posedge lcd_pclk or negedge sys_rst_n)begin
    if(!sys_rst_n)begin
        level_state[0] <= 6'd31;
        level_state[1] <= 6'd32;
    end
    else begin
        if(arrhythmia_level == 2'd0)begin
            level_state[0] <= 6'd31;
            level_state[1] <= 6'd32;
        end
        else begin
            level_state[0] <= 6'd37;
            level_state[1] <= 6'd38;
        end
    end
end

//字体大小位置
localparam CHAR_POS_X  = 11'd322;                 //字符区域起始点横坐标
localparam CHAR_POS_Y  = 11'd43;                 //字符区域起始点纵坐标
localparam CHAR_WIDTH  = 11'd64;               //字符区域宽度
localparam CHAR_HEIGHT = 11'd64;                //字符区域高度

localparam pos_X_remove1  = 11'd104;               //字符区域宽度

// 字符间距参数
localparam CHAR_SPACING = 11'd10;  // 字符间距
localparam CHINESE_WIDTH = 11'd64; // 中文字符宽度64
localparam CHINESE_HEIGHT = 11'd64; // 中文字符高度64
localparam LETTER_WIDTH = 11'd32;  // 英文字母宽度32（修正）
localparam LETTER_HEIGHT = 11'd64; // 英文字母高度64（修正）

// 颜色定义
localparam WHITE  = 24'b11111111_11111111_11111111;  // 白色
localparam BLACK  = 24'b00000000_00000000_00000000;  // 黑色
localparam BLUE   = 24'h0000FF;  // 蓝色
localparam GREEN  = 24'h00FF00;  // 绿色
localparam RED    = 24'hFF0000;  // 红色
localparam GRAY   = 24'h808080;  // 灰色
localparam YELLOW = 24'hFFFF00;  // 黄色
localparam LIGHT_BLUE = 24'hADD8E6; // 浅蓝色
localparam LIGHT_GREEN = 24'h90EE90; // 浅绿色

//主界面色块区域

localparam xinlv_X_START = 11'd56;
localparam xinlv_X_END = 11'd456;
localparam xinlv_Y_START = 11'd175;
localparam xinlv_Y_END = 11'd275;

localparam RR_X_START = 11'd568;
localparam RR_X_END = 11'd968;
localparam RR_Y_START = 11'd175;
localparam RR_Y_END = 11'd275;

localparam HRV_X_START = 11'd56;
localparam HRV_X_END = 11'd456;
localparam HRV_Y_START = 11'd325;
localparam HRV_Y_END = 11'd425;

localparam Level_X_START = 11'd568;
localparam Level_X_END = 11'd968;
localparam Level_Y_START = 11'd325;
localparam Level_Y_END = 11'd425;

localparam xdt_X_START = 11'd62;
localparam xdt_X_END = 11'd412;
localparam xdt_Y_START = 11'd475;
localparam xdt_Y_END = 11'd575;

localparam save_X_START = 11'd487;
localparam save_X_END = 11'd687;
localparam save_Y_START = 11'd475;
localparam save_Y_END = 11'd575;

localparam search_X_START = 11'd762;
localparam search_X_END = 11'd962;
localparam search_Y_START = 11'd475;
localparam search_Y_END = 11'd575;

//子界面色块区域

localparam return_X_START = 11'd72;
localparam return_X_END = 11'd272;
localparam return_Y_START = 11'd25;
localparam return_Y_END = 11'd125;

localparam sel_X_START = 11'd156;
localparam sel_X_END = 11'd356;
localparam sel_Y_START = 11'd495;
localparam sel_Y_END = 11'd595;

localparam del_X_START = 11'd668;
localparam del_X_END = 11'd868;
localparam del_Y_START = 11'd495;
localparam del_Y_END = 11'd595;

localparam data1_X_START = 11'd312;
localparam data1_X_END = 11'd712;
localparam data1_Y_START = 11'd100;
localparam data1_Y_END = 11'd180;

localparam data2_X_START = 11'd312;
localparam data2_X_END = 11'd712;
localparam data2_Y_START = 11'd200;
localparam data2_Y_END = 11'd280;

localparam data3_X_START = 11'd312;
localparam data3_X_END = 11'd712;
localparam data3_Y_START = 11'd300;
localparam data3_Y_END = 11'd380;

localparam data4_X_START = 11'd312;
localparam data4_X_END = 11'd712;
localparam data4_Y_START = 11'd400;
localparam data4_Y_END = 11'd480;

// 文字显示偏移量
localparam TEXT_OFFSET_X = 11'd30;  // 水平偏移
localparam TEXT_OFFSET_Y = 11'd20;  // 垂直偏移

localparam TEXT_OFFSET_X1 = 11'd100;  // 水平偏移
localparam TEXT_OFFSET_Y1 = 11'd5;  // 垂直偏移

// 主界面文字显示位置
localparam XINLV_TEXT_X = xinlv_X_START + TEXT_OFFSET_X;
localparam XINLV_TEXT_Y = xinlv_Y_START + TEXT_OFFSET_Y;

localparam RR_TEXT_X = RR_X_START + TEXT_OFFSET_X;
localparam RR_TEXT_Y = RR_Y_START + TEXT_OFFSET_Y;

localparam HRV_TEXT_X = HRV_X_START + TEXT_OFFSET_X;
localparam HRV_TEXT_Y = HRV_Y_START + TEXT_OFFSET_Y;

localparam LEVEL_TEXT_X = Level_X_START + TEXT_OFFSET_X;
localparam LEVEL_TEXT_Y = Level_Y_START + TEXT_OFFSET_Y;

localparam XDT_TEXT_X = xdt_X_START + TEXT_OFFSET_X;
localparam XDT_TEXT_Y = xdt_Y_START + TEXT_OFFSET_Y;

localparam SAVE_TEXT_X = save_X_START + TEXT_OFFSET_X;
localparam SAVE_TEXT_Y = save_Y_START + TEXT_OFFSET_Y;

localparam SEARCH_TEXT_X = search_X_START + TEXT_OFFSET_X;
localparam SEARCH_TEXT_Y = search_Y_START + TEXT_OFFSET_Y;

// 子界面文字显示位置
localparam RETURN_TEXT_X = return_X_START + TEXT_OFFSET_X;
localparam RETURN_TEXT_Y = return_Y_START + TEXT_OFFSET_Y;

localparam SEL_TEXT_X = sel_X_START + TEXT_OFFSET_X;
localparam SEL_TEXT_Y = sel_Y_START + TEXT_OFFSET_Y;

localparam DEL_TEXT_X = del_X_START + TEXT_OFFSET_X;
localparam DEL_TEXT_Y = del_Y_START + TEXT_OFFSET_Y;

localparam DATA1_TEXT_X = data1_X_START + TEXT_OFFSET_X1;
localparam DATA1_TEXT_Y = data1_Y_START + TEXT_OFFSET_Y1;

localparam DATA2_TEXT_X = data2_X_START + TEXT_OFFSET_X1;
localparam DATA2_TEXT_Y = data2_Y_START + TEXT_OFFSET_Y1;

localparam DATA3_TEXT_X = data3_X_START + TEXT_OFFSET_X1;
localparam DATA3_TEXT_Y = data3_Y_START + TEXT_OFFSET_Y1;

localparam DATA4_TEXT_X = data4_X_START + TEXT_OFFSET_X1;
localparam DATA4_TEXT_Y = data4_Y_START + TEXT_OFFSET_Y1;


reg  [4095:0]  char  [45:0] ;                //字符数组

 //给字符数组赋值，用于存储字模数据
always @(posedge lcd_pclk) begin
    char[0]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h00,
8'h00,8'h1F,8'hF8,8'h00,8'h00,8'h3C,8'h3E,8'h00,8'h00,8'h78,8'h0F,8'h00,8'h00,8'hF0,8'h07,8'h00,
8'h01,8'hE0,8'h07,8'h80,8'h03,8'hE0,8'h03,8'hC0,8'h03,8'hC0,8'h03,8'hC0,8'h07,8'hC0,8'h03,8'hE0,
8'h07,8'hC0,8'h01,8'hE0,8'h07,8'h80,8'h01,8'hE0,8'h0F,8'h80,8'h01,8'hF0,8'h0F,8'h80,8'h01,8'hF0,
8'h0F,8'h80,8'h01,8'hF0,8'h0F,8'h80,8'h00,8'hF0,8'h0F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,
8'h1F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,
8'h1F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,
8'h1F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h00,8'hF8,
8'h1F,8'h00,8'h00,8'hF8,8'h0F,8'h80,8'h00,8'hF0,8'h0F,8'h80,8'h01,8'hF0,8'h0F,8'h80,8'h01,8'hF0,
8'h0F,8'h80,8'h01,8'hF0,8'h07,8'h80,8'h01,8'hE0,8'h07,8'hC0,8'h01,8'hE0,8'h07,8'hC0,8'h03,8'hE0,
8'h03,8'hC0,8'h03,8'hC0,8'h03,8'hE0,8'h03,8'hC0,8'h01,8'hE0,8'h07,8'h80,8'h00,8'hF0,8'h0F,8'h00,
8'h00,8'h78,8'h0E,8'h00,8'h00,8'h3C,8'h3C,8'h00,8'h00,8'h1F,8'hF8,8'h00,8'h00,8'h07,8'hE0,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "0"
    char[1]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h00,
8'h00,8'h00,8'hC0,8'h00,8'h00,8'h01,8'hC0,8'h00,8'h00,8'h07,8'hC0,8'h00,8'h01,8'hFF,8'hC0,8'h00,
8'h01,8'hFF,8'hC0,8'h00,8'h00,8'h07,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h07,8'hE0,8'h00,
8'h00,8'h0F,8'hF0,8'h00,8'h01,8'hFF,8'hFF,8'h80,8'h01,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "1"
    char[2]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hF0,8'h00,
8'h00,8'h3F,8'hFC,8'h00,8'h00,8'hF0,8'h3F,8'h00,8'h01,8'hC0,8'h1F,8'h80,8'h03,8'h80,8'h0F,8'h80,
8'h07,8'h80,8'h07,8'hC0,8'h07,8'h00,8'h07,8'hC0,8'h0F,8'h00,8'h03,8'hE0,8'h0F,8'h00,8'h03,8'hE0,
8'h0F,8'h80,8'h03,8'hE0,8'h0F,8'h80,8'h03,8'hE0,8'h0F,8'hC0,8'h03,8'hE0,8'h0F,8'hC0,8'h03,8'hE0,
8'h0F,8'hC0,8'h03,8'hE0,8'h07,8'h80,8'h03,8'hC0,8'h00,8'h00,8'h07,8'hC0,8'h00,8'h00,8'h07,8'hC0,
8'h00,8'h00,8'h07,8'h80,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h0F,8'h00,8'h00,8'h00,8'h1E,8'h00,
8'h00,8'h00,8'h3C,8'h00,8'h00,8'h00,8'h38,8'h00,8'h00,8'h00,8'h70,8'h00,8'h00,8'h00,8'hE0,8'h00,
8'h00,8'h01,8'hC0,8'h00,8'h00,8'h01,8'hC0,8'h00,8'h00,8'h03,8'h80,8'h00,8'h00,8'h07,8'h00,8'h00,
8'h00,8'h0E,8'h00,8'h00,8'h00,8'h1C,8'h00,8'h00,8'h00,8'h38,8'h00,8'h00,8'h00,8'h70,8'h00,8'h00,
8'h00,8'hE0,8'h00,8'h30,8'h01,8'hC0,8'h00,8'h30,8'h03,8'h80,8'h00,8'h30,8'h03,8'h00,8'h00,8'h30,
8'h07,8'h00,8'h00,8'h60,8'h0E,8'h00,8'h00,8'hE0,8'h0C,8'h00,8'h01,8'hE0,8'h1F,8'hFF,8'hFF,8'hE0,
8'h1F,8'hFF,8'hFF,8'hE0,8'h1F,8'hFF,8'hFF,8'hE0,8'h1F,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "2"
    char[3]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hE0,8'h00,
8'h00,8'h7F,8'hF8,8'h00,8'h00,8'hF0,8'h7C,8'h00,8'h01,8'hC0,8'h3E,8'h00,8'h03,8'h80,8'h1F,8'h00,
8'h03,8'h80,8'h0F,8'h80,8'h07,8'h80,8'h0F,8'h80,8'h07,8'h80,8'h07,8'hC0,8'h07,8'hC0,8'h07,8'hC0,
8'h07,8'hC0,8'h07,8'hC0,8'h07,8'hC0,8'h07,8'hC0,8'h03,8'h80,8'h07,8'hC0,8'h00,8'h00,8'h07,8'hC0,
8'h00,8'h00,8'h07,8'hC0,8'h00,8'h00,8'h07,8'h80,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h0F,8'h00,
8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h3C,8'h00,8'h00,8'h00,8'hF8,8'h00,8'h00,8'h0F,8'hE0,8'h00,
8'h00,8'h0F,8'hF8,8'h00,8'h00,8'h00,8'h7C,8'h00,8'h00,8'h00,8'h1F,8'h00,8'h00,8'h00,8'h0F,8'h80,
8'h00,8'h00,8'h07,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hE0,8'h00,8'h00,8'h01,8'hE0,
8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hF0,
8'h03,8'h80,8'h01,8'hF0,8'h07,8'hC0,8'h01,8'hF0,8'h0F,8'hC0,8'h01,8'hF0,8'h0F,8'hC0,8'h01,8'hE0,
8'h0F,8'hC0,8'h03,8'hE0,8'h0F,8'h80,8'h03,8'hE0,8'h07,8'h80,8'h07,8'hC0,8'h07,8'h80,8'h07,8'h80,
8'h03,8'hC0,8'h0F,8'h00,8'h01,8'hF0,8'h3E,8'h00,8'h00,8'h7F,8'hFC,8'h00,8'h00,8'h1F,8'hE0,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "3"
    char[4]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h0E,8'h00,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h3E,8'h00,
8'h00,8'h00,8'h3E,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,8'hDE,8'h00,8'h00,8'h00,8'hDE,8'h00,
8'h00,8'h01,8'h9E,8'h00,8'h00,8'h03,8'h9E,8'h00,8'h00,8'h03,8'h1E,8'h00,8'h00,8'h06,8'h1E,8'h00,
8'h00,8'h0E,8'h1E,8'h00,8'h00,8'h0C,8'h1E,8'h00,8'h00,8'h18,8'h1E,8'h00,8'h00,8'h18,8'h1E,8'h00,
8'h00,8'h30,8'h1E,8'h00,8'h00,8'h60,8'h1E,8'h00,8'h00,8'h60,8'h1E,8'h00,8'h00,8'hC0,8'h1E,8'h00,
8'h01,8'hC0,8'h1E,8'h00,8'h01,8'h80,8'h1E,8'h00,8'h03,8'h00,8'h1E,8'h00,8'h03,8'h00,8'h1E,8'h00,
8'h06,8'h00,8'h1E,8'h00,8'h0C,8'h00,8'h1E,8'h00,8'h0C,8'h00,8'h1E,8'h00,8'h18,8'h00,8'h1E,8'h00,
8'h3F,8'hFF,8'hFF,8'hFC,8'h3F,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h1E,8'h00,
8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h1E,8'h00,
8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h1E,8'h00,
8'h00,8'h00,8'h3F,8'h00,8'h00,8'h0F,8'hFF,8'hF8,8'h00,8'h0F,8'hFF,8'hF8,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "4"
    char[5]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h01,8'hFF,8'hFF,8'hE0,8'h01,8'hFF,8'hFF,8'hE0,8'h01,8'hFF,8'hFF,8'hE0,8'h01,8'hFF,8'hFF,8'hC0,
8'h01,8'h80,8'h00,8'h00,8'h01,8'h80,8'h00,8'h00,8'h01,8'h80,8'h00,8'h00,8'h01,8'h80,8'h00,8'h00,
8'h01,8'h80,8'h00,8'h00,8'h01,8'h80,8'h00,8'h00,8'h01,8'h80,8'h00,8'h00,8'h01,8'h80,8'h00,8'h00,
8'h03,8'h00,8'h00,8'h00,8'h03,8'h00,8'h00,8'h00,8'h03,8'h00,8'h00,8'h00,8'h03,8'h00,8'h00,8'h00,
8'h03,8'h03,8'hF8,8'h00,8'h03,8'h1F,8'hFE,8'h00,8'h03,8'h3F,8'hFF,8'h00,8'h03,8'h78,8'h1F,8'h80,
8'h03,8'hE0,8'h0F,8'hC0,8'h03,8'hC0,8'h07,8'hC0,8'h03,8'h80,8'h03,8'hE0,8'h03,8'h00,8'h03,8'hE0,
8'h00,8'h00,8'h03,8'hE0,8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hF0,
8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hF0,8'h03,8'h80,8'h01,8'hF0,
8'h07,8'hC0,8'h01,8'hF0,8'h0F,8'hC0,8'h01,8'hF0,8'h0F,8'hC0,8'h01,8'hE0,8'h0F,8'hC0,8'h03,8'hE0,
8'h0F,8'h80,8'h03,8'hE0,8'h0F,8'h80,8'h03,8'hC0,8'h07,8'h80,8'h07,8'hC0,8'h03,8'h80,8'h07,8'h80,
8'h01,8'hC0,8'h0F,8'h00,8'h00,8'hF0,8'h3E,8'h00,8'h00,8'h7F,8'hFC,8'h00,8'h00,8'h0F,8'hF0,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "5"
    char[6]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'hFC,8'h00,
8'h00,8'h07,8'hFF,8'h00,8'h00,8'h1F,8'h07,8'h80,8'h00,8'h3C,8'h03,8'hC0,8'h00,8'h70,8'h03,8'hE0,
8'h00,8'hE0,8'h03,8'hE0,8'h01,8'hE0,8'h03,8'hE0,8'h01,8'hC0,8'h03,8'hE0,8'h03,8'hC0,8'h01,8'hC0,
8'h03,8'h80,8'h00,8'h00,8'h07,8'h80,8'h00,8'h00,8'h07,8'h80,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,
8'h0F,8'h80,8'h00,8'h00,8'h0F,8'h00,8'h00,8'h00,8'h0F,8'h00,8'h00,8'h00,8'h0F,8'h01,8'hF8,8'h00,
8'h1F,8'h0F,8'hFF,8'h00,8'h1F,8'h1F,8'hFF,8'h80,8'h1F,8'h3E,8'h0F,8'hC0,8'h1F,8'h78,8'h03,8'hE0,
8'h1F,8'h60,8'h01,8'hE0,8'h1F,8'hC0,8'h01,8'hF0,8'h1F,8'hC0,8'h00,8'hF0,8'h1F,8'h80,8'h00,8'hF0,
8'h1F,8'h80,8'h00,8'h78,8'h1F,8'h00,8'h00,8'h78,8'h1F,8'h00,8'h00,8'h78,8'h1F,8'h00,8'h00,8'h78,
8'h1F,8'h00,8'h00,8'h78,8'h1F,8'h00,8'h00,8'h78,8'h0F,8'h00,8'h00,8'h78,8'h0F,8'h00,8'h00,8'h78,
8'h0F,8'h80,8'h00,8'h78,8'h0F,8'h80,8'h00,8'h78,8'h07,8'h80,8'h00,8'h70,8'h07,8'hC0,8'h00,8'hF0,
8'h07,8'hC0,8'h00,8'hF0,8'h03,8'hE0,8'h00,8'hE0,8'h03,8'hE0,8'h01,8'hE0,8'h01,8'hF0,8'h01,8'hC0,
8'h00,8'hF8,8'h03,8'h80,8'h00,8'h7E,8'h0F,8'h00,8'h00,8'h1F,8'hFC,8'h00,8'h00,8'h07,8'hF0,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "6"
    char[7]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h03,8'hFF,8'hFF,8'hF0,8'h07,8'hFF,8'hFF,8'hF0,8'h07,8'hFF,8'hFF,8'hF0,8'h07,8'hFF,8'hFF,8'hE0,
8'h07,8'h80,8'h00,8'hC0,8'h07,8'h00,8'h00,8'hC0,8'h06,8'h00,8'h01,8'h80,8'h06,8'h00,8'h01,8'h80,
8'h0C,8'h00,8'h03,8'h00,8'h0C,8'h00,8'h03,8'h00,8'h0C,8'h00,8'h06,8'h00,8'h00,8'h00,8'h06,8'h00,
8'h00,8'h00,8'h0C,8'h00,8'h00,8'h00,8'h1C,8'h00,8'h00,8'h00,8'h18,8'h00,8'h00,8'h00,8'h38,8'h00,
8'h00,8'h00,8'h38,8'h00,8'h00,8'h00,8'h30,8'h00,8'h00,8'h00,8'h70,8'h00,8'h00,8'h00,8'h70,8'h00,
8'h00,8'h00,8'hE0,8'h00,8'h00,8'h00,8'hE0,8'h00,8'h00,8'h01,8'hE0,8'h00,8'h00,8'h01,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'h80,8'h00,8'h00,8'h07,8'h80,8'h00,
8'h00,8'h07,8'h80,8'h00,8'h00,8'h07,8'h80,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h0F,8'h80,8'h00,
8'h00,8'h0F,8'h80,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h1F,8'h80,8'h00,
8'h00,8'h1F,8'h80,8'h00,8'h00,8'h1F,8'h80,8'h00,8'h00,8'h1F,8'h80,8'h00,8'h00,8'h1F,8'h80,8'h00,
8'h00,8'h1F,8'h80,8'h00,8'h00,8'h1F,8'h80,8'h00,8'h00,8'h1F,8'h80,8'h00,8'h00,8'h0F,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "7"
    char[8]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hF0,8'h00,
8'h00,8'h7F,8'hFE,8'h00,8'h00,8'hF8,8'h1F,8'h00,8'h01,8'hE0,8'h07,8'h80,8'h03,8'hC0,8'h03,8'hC0,
8'h07,8'h80,8'h01,8'hE0,8'h07,8'h80,8'h01,8'hE0,8'h0F,8'h00,8'h00,8'hF0,8'h0F,8'h00,8'h00,8'hF0,
8'h0F,8'h00,8'h00,8'hF0,8'h0F,8'h00,8'h00,8'hF0,8'h0F,8'h00,8'h00,8'hF0,8'h0F,8'h80,8'h00,8'hF0,
8'h0F,8'h80,8'h00,8'hF0,8'h07,8'hC0,8'h01,8'hE0,8'h07,8'hE0,8'h01,8'hE0,8'h03,8'hF0,8'h01,8'hC0,
8'h01,8'hFC,8'h03,8'h80,8'h00,8'hFE,8'h07,8'h00,8'h00,8'h7F,8'hCE,8'h00,8'h00,8'h3F,8'hFC,8'h00,
8'h00,8'h1F,8'hF8,8'h00,8'h00,8'h73,8'hFE,8'h00,8'h00,8'hE0,8'hFF,8'h00,8'h01,8'hC0,8'h3F,8'h80,
8'h03,8'hC0,8'h1F,8'hC0,8'h07,8'h80,8'h07,8'hE0,8'h07,8'h00,8'h03,8'hE0,8'h0F,8'h00,8'h01,8'hF0,
8'h0F,8'h00,8'h01,8'hF0,8'h1E,8'h00,8'h00,8'hF8,8'h1E,8'h00,8'h00,8'h78,8'h1E,8'h00,8'h00,8'h78,
8'h1E,8'h00,8'h00,8'h78,8'h1E,8'h00,8'h00,8'h78,8'h1E,8'h00,8'h00,8'h78,8'h1E,8'h00,8'h00,8'h78,
8'h0F,8'h00,8'h00,8'h70,8'h0F,8'h00,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hE0,8'h03,8'hC0,8'h01,8'hE0,
8'h01,8'hE0,8'h03,8'hC0,8'h00,8'hF8,8'h0F,8'h00,8'h00,8'h3F,8'hFE,8'h00,8'h00,8'h0F,8'hF0,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "8"
    char[9]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hE0,8'h00,
8'h00,8'h7F,8'hFC,8'h00,8'h00,8'hF0,8'h3E,8'h00,8'h01,8'hE0,8'h0F,8'h00,8'h03,8'hC0,8'h07,8'h80,
8'h07,8'h80,8'h03,8'hC0,8'h07,8'h00,8'h03,8'hC0,8'h0F,8'h00,8'h01,8'hE0,8'h0F,8'h00,8'h01,8'hE0,
8'h0E,8'h00,8'h01,8'hF0,8'h1E,8'h00,8'h00,8'hF0,8'h1E,8'h00,8'h00,8'hF0,8'h1E,8'h00,8'h00,8'hF0,
8'h1E,8'h00,8'h00,8'hF8,8'h1E,8'h00,8'h00,8'hF8,8'h1E,8'h00,8'h00,8'hF8,8'h1E,8'h00,8'h00,8'hF8,
8'h1E,8'h00,8'h00,8'hF8,8'h1E,8'h00,8'h01,8'hF8,8'h1F,8'h00,8'h01,8'hF8,8'h0F,8'h00,8'h03,8'hF8,
8'h0F,8'h80,8'h07,8'hF8,8'h0F,8'h80,8'h0E,8'hF8,8'h07,8'hC0,8'h1E,8'hF8,8'h03,8'hF0,8'h7C,8'hF8,
8'h01,8'hFF,8'hF8,8'hF8,8'h00,8'hFF,8'hE0,8'hF8,8'h00,8'h3F,8'h81,8'hF0,8'h00,8'h00,8'h01,8'hF0,
8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h01,8'hE0,
8'h00,8'h00,8'h03,8'hE0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h03,8'h80,8'h07,8'hC0,
8'h07,8'hC0,8'h07,8'h80,8'h07,8'hC0,8'h0F,8'h00,8'h07,8'hC0,8'h0F,8'h00,8'h07,8'hC0,8'h1E,8'h00,
8'h03,8'hC0,8'h3C,8'h00,8'h03,8'hE0,8'hF8,8'h00,8'h00,8'hFF,8'hE0,8'h00,8'h00,8'h3F,8'h80,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "9"
    char[10]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hF0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h01,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'hFC,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h01,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hFC,8'h07,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h03,8'hF8,8'h0F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h03,8'hF8,8'h0F,8'hE0,8'h00,
8'h00,8'h00,8'h00,8'h07,8'hF0,8'h1F,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h1F,8'hE0,8'h00,
8'h00,8'h60,8'hE0,8'h07,8'hE0,8'h1F,8'hC0,8'h00,8'h00,8'h61,8'hF0,8'h0F,8'hC0,8'h3F,8'hC0,8'h00,
8'h00,8'h61,8'hF0,8'h0F,8'h80,8'h3F,8'h80,8'h00,8'h00,8'hE1,8'hF8,8'h1F,8'h00,8'h7F,8'h00,8'h00,
8'h00,8'hE1,8'hF8,8'h3E,8'h00,8'h7F,8'h00,8'h00,8'h01,8'hE1,8'hFC,8'h7C,8'h00,8'hFE,8'h00,8'h00,
8'h01,8'hE1,8'hFE,8'hF8,8'h01,8'hFC,8'h00,8'h00,8'h03,8'hE3,8'hFF,8'hE0,8'h01,8'hF8,8'h00,8'h00,
8'h03,8'hE1,8'hFF,8'hC0,8'h03,8'hF0,8'h00,8'h00,8'h07,8'hE0,8'h0F,8'hF0,8'h07,8'hE0,8'h00,8'h00,
8'h07,8'hE0,8'h03,8'hFC,8'h0F,8'h80,8'h00,8'h00,8'h0F,8'hE0,8'h01,8'hFE,8'h0F,8'h00,8'h00,8'h00,
8'h0F,8'hE0,8'h00,8'h7F,8'h9E,8'h00,8'h00,8'h00,8'h1F,8'hE0,8'h00,8'h3F,8'hFC,8'h00,8'h00,8'h00,
8'h1F,8'hC0,8'h00,8'h1F,8'hFE,8'h00,8'h00,8'h00,8'h3F,8'hC0,8'h00,8'h0F,8'hFF,8'hC0,8'h00,8'h0E,
8'h3F,8'hC0,8'h00,8'h03,8'hFF,8'hFF,8'h01,8'hFC,8'h3F,8'h80,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFC,
8'h3F,8'h80,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'hFC,8'h3F,8'h00,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'hF8,
8'h3E,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hF8,8'h18,8'h00,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hF0,
8'h00,8'h00,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hE0,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hFE,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h70,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "心"
    char[11]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h01,8'hC0,8'h1C,8'h00,8'h00,8'h00,8'h00,8'h01,8'h03,8'hE0,8'h3E,8'h00,8'h00,8'h00,
8'h00,8'h03,8'h87,8'hE0,8'h3E,8'h00,8'h00,8'h00,8'h00,8'h07,8'hC3,8'hE0,8'h7E,8'h00,8'h00,8'h00,
8'h00,8'h07,8'hC3,8'hE0,8'h7F,8'hFF,8'hF8,8'h00,8'h00,8'h07,8'hC3,8'hE0,8'hFF,8'hFF,8'hF8,8'h00,
8'h00,8'h07,8'hC3,8'hE1,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h07,8'hC3,8'hE3,8'hE0,8'h00,8'h00,8'h00,
8'h00,8'h07,8'hC3,8'hE7,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h07,8'hC3,8'hEF,8'h00,8'hE0,8'h00,8'h00,
8'h00,8'h03,8'hC3,8'hE4,8'hC1,8'hF8,8'h00,8'h00,8'h00,8'h03,8'hC3,8'hE1,8'hE1,8'hFC,8'h00,8'h00,
8'h00,8'h03,8'hC3,8'hC7,8'hE0,8'h7F,8'h00,8'h00,8'h00,8'h03,8'hC3,8'h8F,8'hC0,8'h0F,8'h00,8'h00,
8'h00,8'h03,8'h80,8'h3F,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h03,8'h00,8'hFF,8'hFC,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h07,8'hF1,8'hFF,8'h80,8'h00,8'h00,8'h00,8'h00,8'h1F,8'hC0,8'h3F,8'hF0,8'h00,8'h00,
8'h00,8'h00,8'hFF,8'h80,8'h07,8'hFE,8'h00,8'h00,8'h00,8'h07,8'hFE,8'h00,8'h00,8'hFF,8'hF0,8'h00,
8'h00,8'h7F,8'hFB,8'hFF,8'hFF,8'h3F,8'hFF,8'hC0,8'h0F,8'hFF,8'hE3,8'hFF,8'hFF,8'h8F,8'hFF,8'hFC,
8'h1F,8'hFF,8'h83,8'hFF,8'hFC,8'h01,8'hFF,8'hFC,8'h1F,8'hFE,8'h00,8'h0F,8'hE0,8'h00,8'h7F,8'hF8,
8'h0F,8'hF0,8'h40,8'h0F,8'hE0,8'h00,8'h1F,8'hF0,8'h07,8'hC0,8'hFF,8'hFF,8'hFF,8'hF8,8'h07,8'hF0,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFE,8'h03,8'hE0,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h38,8'h0F,8'hE0,8'h38,8'h00,8'h00,
8'h00,8'h00,8'h3E,8'h0F,8'hE0,8'h78,8'h00,8'h00,8'h00,8'h00,8'h3F,8'h0F,8'hE1,8'hF8,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'hCF,8'hE3,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hCF,8'hE7,8'hC0,8'h00,8'h00,
8'h00,8'h07,8'h80,8'h0F,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,8'h00,
8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,
8'h00,8'h1F,8'h00,8'h00,8'h00,8'h1F,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "鉴"
    char[12]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h01,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,
8'h00,8'h00,8'h04,8'h00,8'h03,8'hF8,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'h00,8'h03,8'hF8,8'h00,8'h00,
8'h07,8'hFF,8'hFF,8'h80,8'h03,8'hF8,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'h80,8'h01,8'hF8,8'h00,8'h00,
8'h0F,8'hFF,8'hFF,8'h80,8'h01,8'hF8,8'h00,8'h00,8'h0E,8'h00,8'h3F,8'h81,8'h01,8'hF8,8'h08,8'h00,
8'h00,8'h20,8'h1F,8'h87,8'hFF,8'hFF,8'hFE,8'h00,8'h00,8'hF8,8'h1F,8'h0F,8'hFF,8'hFF,8'hFF,8'h00,
8'h00,8'hF8,8'h1F,8'h0F,8'hFF,8'hFF,8'hFF,8'h00,8'h01,8'hF8,8'h1F,8'h0F,8'hFF,8'hFF,8'hFF,8'h00,
8'h01,8'hF8,8'h1F,8'h0F,8'hC0,8'hF0,8'h7F,8'h00,8'h01,8'hF8,8'h1F,8'h07,8'hC0,8'hF0,8'h3E,8'h00,
8'h01,8'hF8,8'h1F,8'h07,8'hC0,8'hF0,8'h3E,8'h00,8'h01,8'hF0,8'h1E,8'h07,8'hC0,8'hF0,8'h3E,8'h00,
8'h01,8'hF0,8'h1E,8'h07,8'hC1,8'hF0,8'h3E,8'h00,8'h01,8'hF0,8'h1E,8'h07,8'hE1,8'hF0,8'h7E,8'h00,
8'h01,8'hF0,8'h1E,8'h07,8'hFF,8'hFF,8'hFE,8'h00,8'h01,8'hF0,8'h1E,8'h07,8'hFF,8'hFF,8'hFE,8'h00,
8'h03,8'hFF,8'hFF,8'hE7,8'hFF,8'hFF,8'hFE,8'h00,8'h03,8'hFF,8'hFF,8'hF3,8'hE1,8'hFF,8'hFC,8'h00,
8'h03,8'hFF,8'hFF,8'hF1,8'h01,8'hE0,8'h18,8'h00,8'h03,8'hF8,8'h1F,8'hF0,8'hF3,8'hE0,8'h00,8'h00,
8'h00,8'hC0,8'h03,8'hF1,8'hFB,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h01,8'hF0,8'h7F,8'hC0,8'h00,8'h00,
8'h00,8'h00,8'h01,8'hF0,8'h3F,8'hC0,8'h00,8'h00,8'h1F,8'hFF,8'hF9,8'hF0,8'h0F,8'hE0,8'h00,8'h00,
8'h3F,8'hFF,8'hF9,8'hE0,8'h0F,8'hF8,8'h00,8'h00,8'h3F,8'hFF,8'hC3,8'hE0,8'h1F,8'hFE,8'h00,8'h00,
8'h7F,8'hFE,8'h03,8'hE0,8'h1F,8'hFF,8'h80,8'h00,8'h3F,8'hE0,8'h03,8'hE0,8'h3F,8'h7F,8'hE0,8'h00,
8'h1E,8'h00,8'h07,8'hC0,8'h7E,8'h3F,8'hFC,8'h00,8'h00,8'h00,8'h0F,8'hC1,8'hFC,8'h0F,8'hFF,8'hF0,
8'h00,8'h20,8'h1F,8'hC3,8'hF8,8'h07,8'hFF,8'hFC,8'h00,8'h1F,8'hFF,8'h9F,8'hF0,8'h03,8'hFF,8'hFC,
8'h00,8'h1F,8'hFF,8'hBF,8'hE0,8'h00,8'hFF,8'hF8,8'h00,8'h0F,8'hFF,8'h1F,8'h80,8'h00,8'h7F,8'hF0,
8'h00,8'h07,8'hFE,8'h04,8'h00,8'h00,8'h3F,8'hE0,8'h00,8'h00,8'h70,8'h00,8'h00,8'h00,8'h0F,8'hC0,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "驶"
    char[13]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h08,8'h00,8'h00,8'h3F,8'h80,8'h00,8'h00,
8'h00,8'h3E,8'h00,8'h00,8'h7F,8'hE0,8'h00,8'h00,8'h00,8'h7F,8'h00,8'h00,8'hFF,8'hF8,8'h00,8'h00,
8'h00,8'h7F,8'hC0,8'h01,8'hFF,8'hFE,8'h00,8'h00,8'h00,8'h7F,8'hE0,8'h03,8'hF0,8'h7F,8'h80,8'h00,
8'h00,8'h3F,8'hF0,8'h0F,8'hE0,8'h1F,8'hE0,8'h00,8'h00,8'h07,8'hFC,8'h1F,8'h80,8'h07,8'hF8,8'h00,
8'h00,8'h00,8'h40,8'h3F,8'h00,8'h01,8'hFE,8'h00,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hF8,8'h7F,8'h00,
8'h00,8'h00,8'h03,8'hF7,8'hFF,8'hFE,8'h1F,8'h80,8'h00,8'h00,8'h07,8'hE7,8'hFF,8'hFC,8'h03,8'h80,
8'h01,8'hE0,8'hE1,8'h02,8'h1F,8'h80,8'h00,8'h00,8'h07,8'hFF,8'hF0,8'h00,8'h1F,8'h80,8'h00,8'h00,
8'h0F,8'hFF,8'hF8,8'h00,8'h1F,8'hC0,8'h00,8'h00,8'h0F,8'hFF,8'hF8,8'h3F,8'hFF,8'hFF,8'hE0,8'h00,
8'h0F,8'h81,8'hF8,8'h3F,8'hFF,8'hFF,8'hF0,8'h00,8'h0E,8'h01,8'hE0,8'h7F,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h1F,8'h80,8'h00,8'h00,8'h00,8'h07,8'hC0,8'h06,8'h1F,8'h80,8'h00,8'h00,
8'h00,8'h07,8'h80,8'h07,8'h9F,8'h87,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h0F,8'h1F,8'h8F,8'h80,8'h00,
8'h00,8'h07,8'hC0,8'h1F,8'h1F,8'h8F,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h3E,8'h1F,8'h8F,8'hF0,8'h00,
8'h00,8'h01,8'hC0,8'h7C,8'h0F,8'h87,8'hF8,8'h00,8'h00,8'h01,8'h81,8'hF3,8'hBF,8'h83,8'hFC,8'h00,
8'h00,8'h03,8'h83,8'hC1,8'hFF,8'h80,8'hFE,8'h00,8'h07,8'hFF,8'hE0,8'h00,8'hFF,8'h80,8'h1E,8'h00,
8'h1F,8'hFF,8'hFF,8'h00,8'h1F,8'h80,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'hFE,8'h02,8'h00,8'h00,8'h00,
8'h3F,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h00,8'h3F,8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'h80,8'h00,
8'h3C,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFC,8'h30,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'hF8,
8'h00,8'h00,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hE0,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFF,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "途"
    char[14]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h38,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'h00,8'hFC,8'h00,8'h1E,8'h00,8'h00,
8'h01,8'hFE,8'h00,8'hFC,8'h03,8'hFF,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,
8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,
8'h07,8'hFF,8'hFF,8'hFC,8'h00,8'h3F,8'h80,8'h00,8'h03,8'hF8,8'h00,8'hF8,8'h00,8'h1F,8'h80,8'h00,
8'h03,8'hF8,8'h00,8'hF8,8'h00,8'h1F,8'h80,8'h00,8'h03,8'hF8,8'h00,8'hF8,8'h00,8'h1F,8'h80,8'h00,
8'h01,8'hF8,8'h01,8'hFC,8'h00,8'h1F,8'h80,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,
8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,
8'h01,8'hF8,8'h00,8'hF8,8'h00,8'h1F,8'h00,8'h00,8'h00,8'hF8,8'h00,8'hF8,8'h00,8'h1F,8'h00,8'h00,
8'h00,8'hF8,8'h00,8'hF8,8'h00,8'h1F,8'h00,8'h00,8'h00,8'hF8,8'h00,8'hF8,8'h00,8'h3F,8'h00,8'h00,
8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,
8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,8'h00,
8'h00,8'h7F,8'hFF,8'hFC,8'h01,8'hFC,8'h00,8'h00,8'h00,8'h7F,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h38,8'h00,8'hFE,8'h00,8'h00,8'h00,8'h04,8'h00,8'h00,8'h00,8'hFE,8'h00,8'h00,8'h00,8'h0C,
8'h00,8'h00,8'h00,8'h7F,8'hC0,8'h00,8'h00,8'h78,8'h00,8'h00,8'h00,8'h7F,8'hF0,8'h00,8'h03,8'hF8,
8'h00,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hF0,
8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hE0,
8'h00,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'h80,
8'h00,8'h00,8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'hFF,8'hFC,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "电"
    char[15]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1F,8'hC0,8'h00,8'h00,
8'h00,8'h7C,8'h00,8'h00,8'h1F,8'hC0,8'h00,8'h00,8'h00,8'hFE,8'h00,8'hE0,8'h1F,8'hC0,8'h00,8'h00,
8'h00,8'hFF,8'h01,8'hF1,8'hFF,8'hF8,8'h00,8'h00,8'h00,8'hFF,8'hC1,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,
8'h00,8'h7F,8'hE0,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,8'h00,8'h3F,8'hF8,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,
8'h00,8'h0F,8'hFC,8'hF8,8'h0F,8'h80,8'h3E,8'h00,8'h00,8'h00,8'h10,8'hF8,8'h0F,8'h80,8'h1E,8'h00,
8'h00,8'h00,8'h00,8'hF8,8'h0F,8'h80,8'h1E,8'h00,8'h0C,8'h00,8'h00,8'hF8,8'h0F,8'h80,8'h1E,8'h00,
8'h1F,8'h80,8'h00,8'hF8,8'h0F,8'h80,8'h1E,8'h00,8'h1F,8'hE0,8'h00,8'hF8,8'h0F,8'h80,8'h1E,8'h00,
8'h1F,8'hF8,8'h00,8'hF9,8'h0F,8'hFE,8'h1C,8'h00,8'h1F,8'hFC,8'h00,8'hF3,8'hFF,8'hFF,8'h1C,8'h00,
8'h1F,8'hFF,8'h00,8'hF3,8'hFF,8'hFF,8'h80,8'h00,8'h1F,8'hFF,8'h80,8'hF7,8'hF8,8'h3F,8'h80,8'h00,
8'h07,8'hFF,8'hE0,8'hF1,8'hC0,8'h1F,8'h80,8'h00,8'h01,8'hFF,8'h00,8'hF3,8'hE0,8'h1F,8'h80,8'h00,
8'h00,8'h00,8'h00,8'hF3,8'hF0,8'h3F,8'h00,8'h00,8'h00,8'h00,8'h00,8'hF0,8'hF8,8'h3E,8'h00,8'h00,
8'h00,8'h00,8'h01,8'hE0,8'h7C,8'h7E,8'h00,8'h00,8'h00,8'h00,8'h61,8'hE0,8'h1F,8'hFC,8'h00,8'h00,
8'h00,8'h01,8'hE3,8'hE0,8'h0F,8'hF8,8'h00,8'h00,8'h00,8'h0F,8'hE3,8'hE0,8'h07,8'hF8,8'h00,8'h00,
8'h00,8'h3F,8'hC7,8'hC0,8'h03,8'hFC,8'h00,8'h00,8'h01,8'hFF,8'h87,8'hC0,8'h07,8'hFF,8'h00,8'h00,
8'h07,8'hFF,8'h0F,8'h80,8'h0F,8'hFF,8'hC0,8'h00,8'h0F,8'hFE,8'h1F,8'h80,8'h1F,8'hFF,8'hF0,8'h00,
8'h0F,8'hFC,8'h3F,8'h00,8'h3F,8'h3F,8'hFC,8'h00,8'h0F,8'hF0,8'h7E,8'h00,8'hFE,8'h1F,8'hFF,8'hC0,
8'h07,8'hC1,8'hFE,8'h03,8'hFC,8'h0F,8'hFF,8'hFE,8'h00,8'h01,8'hF8,8'h1F,8'hF8,8'h07,8'hFF,8'hFC,
8'h00,8'h00,8'h00,8'h7F,8'hF0,8'h01,8'hFF,8'hF8,8'h00,8'h00,8'h00,8'h7F,8'hC0,8'h00,8'hFF,8'hF0,
8'h00,8'h00,8'h00,8'h3F,8'h00,8'h00,8'h7F,8'hF0,8'h00,8'h00,8'h00,8'h08,8'h00,8'h00,8'h1F,8'hE0,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "波"
    char[16]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'hF0,8'h00,8'h7F,8'h80,
8'h00,8'h7F,8'hFF,8'hFF,8'hF8,8'h01,8'hFF,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hF8,8'h07,8'hFE,8'h00,
8'h00,8'hFF,8'hFF,8'hFF,8'hF0,8'h1F,8'hFC,8'h00,8'h00,8'h01,8'hE0,8'h7C,8'h00,8'hFF,8'hE0,8'h00,
8'h00,8'h01,8'hE0,8'h7C,8'h07,8'hFF,8'h80,8'h00,8'h00,8'h01,8'hE0,8'h7C,8'h0F,8'hFC,8'h00,8'h00,
8'h00,8'h01,8'hE0,8'h7C,8'h07,8'hE0,8'h00,8'h00,8'h00,8'h01,8'hE0,8'h7C,8'h00,8'h00,8'h06,8'h00,
8'h00,8'h01,8'hE0,8'h7C,8'h00,8'h00,8'h1F,8'h00,8'h00,8'h01,8'hE0,8'h7C,8'h00,8'h00,8'h3F,8'h00,
8'h07,8'h03,8'hFF,8'hFF,8'hF8,8'h00,8'h7F,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'hFF,8'h00,
8'h1F,8'hFF,8'hFF,8'hFF,8'hFC,8'h03,8'hFC,8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hF8,8'h0F,8'hF8,8'h00,
8'h3F,8'hFF,8'hFF,8'hFC,8'h00,8'h1F,8'hE0,8'h00,8'h00,8'h03,8'hE0,8'h7C,8'h00,8'h7F,8'h80,8'h78,
8'h00,8'h03,8'hE0,8'h7C,8'h03,8'hFE,8'h00,8'h78,8'h00,8'h03,8'hE0,8'h7C,8'h0F,8'hF8,8'h00,8'hFC,
8'h00,8'h03,8'hE0,8'h7C,8'h0F,8'hC0,8'h01,8'hFC,8'h00,8'h03,8'hE0,8'h7C,8'h02,8'h00,8'h03,8'hF8,
8'h00,8'h07,8'hE0,8'h7C,8'h00,8'h00,8'h07,8'hF8,8'h00,8'h07,8'hC0,8'h7C,8'h00,8'h00,8'h0F,8'hF0,
8'h00,8'h0F,8'hC0,8'h7C,8'h00,8'h00,8'h1F,8'hC0,8'h00,8'h0F,8'hC0,8'h7C,8'h00,8'h00,8'h7F,8'h80,
8'h00,8'h1F,8'hC0,8'h7C,8'h00,8'h00,8'hFF,8'h00,8'h00,8'h3F,8'h80,8'h7C,8'h00,8'h03,8'hFE,8'h00,
8'h00,8'hFF,8'h00,8'h7C,8'h00,8'h0F,8'hF8,8'h00,8'h07,8'hFF,8'h00,8'h7C,8'h00,8'h7F,8'hF0,8'h00,
8'h3F,8'hFE,8'h00,8'h7C,8'h01,8'hFF,8'hE0,8'h00,8'h3F,8'hFC,8'h00,8'h7C,8'h1F,8'hFF,8'h80,8'h00,
8'h1F,8'hF0,8'h00,8'h7C,8'hFF,8'hFE,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h7C,8'hFF,8'hF8,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h78,8'h3F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "形"
    char[17]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h0C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1E,8'h00,8'h04,8'h00,8'h00,8'h20,8'h00,
8'h00,8'h3F,8'h00,8'h0F,8'hFF,8'hFF,8'hF8,8'h00,8'h00,8'h3F,8'hC0,8'h1F,8'hFF,8'hFF,8'hF8,8'h00,
8'h00,8'h3F,8'hE0,8'h3F,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h1F,8'hF8,8'h7F,8'hE0,8'h01,8'hFC,8'h00,
8'h00,8'h07,8'hFC,8'h38,8'h00,8'h00,8'hF8,8'h00,8'h00,8'h00,8'hF8,8'h30,8'h00,8'h00,8'hF8,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hF0,8'h00,
8'h00,8'h02,8'h00,8'h00,8'h00,8'h00,8'hF0,8'h00,8'h00,8'h07,8'hC0,8'h03,8'hC0,8'h00,8'hF0,8'h00,
8'h1F,8'hFF,8'hE0,8'h03,8'hE0,8'h01,8'hF0,8'h00,8'h1F,8'hFF,8'hE0,8'h07,8'hFF,8'hFF,8'hF8,8'h00,
8'h3F,8'hFF,8'hE0,8'h07,8'hFF,8'hFF,8'hF0,8'h00,8'h3E,8'h3F,8'hC0,8'h07,8'hF0,8'h1F,8'hF0,8'h00,
8'h38,8'h0F,8'h80,8'h07,8'h80,8'h00,8'hE0,8'h00,8'h00,8'h0F,8'h80,8'h0F,8'h80,8'h00,8'h00,8'h00,
8'h00,8'h0F,8'h80,8'h0F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h0F,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h0F,8'h80,8'h0F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h0E,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h0F,8'h80,8'h0E,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'hCF,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h0F,8'h81,8'hCF,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h83,8'h8F,8'h80,8'h00,8'h00,8'h0C,
8'h00,8'h0F,8'h87,8'h8F,8'hC0,8'h00,8'h00,8'h3C,8'h00,8'h0F,8'h9F,8'h0F,8'hF0,8'h00,8'h00,8'h7C,
8'h00,8'h0F,8'hFE,8'h07,8'hFE,8'h00,8'h01,8'hFC,8'h00,8'h1F,8'hFC,8'h03,8'hFF,8'hF0,8'h07,8'hFC,
8'h00,8'h3F,8'hFC,8'h01,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'h7F,8'hF8,8'h00,8'h7F,8'hFF,8'hFF,8'hF8,
8'h00,8'h7F,8'hF0,8'h00,8'h3F,8'hFF,8'hFF,8'hF8,8'h00,8'h7F,8'hE0,8'h00,8'h0F,8'hFF,8'hFF,8'hF0,
8'h00,8'h3F,8'hC0,8'h00,8'h03,8'hFF,8'hFF,8'hF0,8'h00,8'h3F,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hE0,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFE,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "记"
    char[18]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h00,8'h00,8'h38,8'h00,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,8'h00,8'h00,8'h03,8'hE0,8'h00,8'h01,8'hFE,8'h00,8'h00,
8'h00,8'h01,8'h80,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h00,8'h00,8'hFF,8'hE0,8'h00,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'hC0,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,
8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,
8'h3F,8'hFF,8'hC0,8'h0F,8'hFF,8'hFF,8'hFF,8'hF8,8'h3F,8'hC0,8'h00,8'h0F,8'hE0,8'h0F,8'hFF,8'hE0,
8'h3C,8'h00,8'hC0,8'h0F,8'hE0,8'h38,8'h7F,8'hC0,8'h00,8'h01,8'hF0,8'h0F,8'hE0,8'h3C,8'h06,8'h00,
8'h00,8'h03,8'hF8,8'h0F,8'hE0,8'h7C,8'h00,8'h00,8'h00,8'h01,8'hFE,8'h0F,8'hE0,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'hFF,8'h8F,8'hF1,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h3F,8'hFB,8'hE0,8'h00,8'h00,
8'h00,8'h00,8'h00,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'h80,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'hEF,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'h00,8'hFF,8'h8F,8'hE7,8'hF0,8'h00,8'h00,
8'h00,8'h3F,8'hFF,8'h0F,8'hE1,8'hF8,8'h00,8'h00,8'h00,8'h7F,8'hFC,8'h0F,8'hE0,8'hFE,8'h00,8'h00,
8'h00,8'hFF,8'hF0,8'h0F,8'hE0,8'h3F,8'h00,8'h00,8'h00,8'hFF,8'hC0,8'h0F,8'hE0,8'h0F,8'hC0,8'h00,
8'h00,8'hFF,8'h00,8'h0F,8'hE0,8'h03,8'hE0,8'h00,8'h00,8'hFC,8'h00,8'h0F,8'hE0,8'h01,8'hF8,8'h00,
8'h00,8'h00,8'h0F,8'h3F,8'hE0,8'h00,8'h78,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h07,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hFF,8'h80,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "录"
    char[19]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h07,8'h80,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h07,8'hC0,8'h00,8'h00,
8'h00,8'h07,8'hE0,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h0F,8'hE0,8'h00,8'h00,
8'h00,8'h07,8'hE0,8'h00,8'h1F,8'hC0,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h1F,8'hC0,8'h00,8'h00,
8'h00,8'h07,8'hE0,8'h00,8'h3F,8'h80,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h7F,8'h80,8'h00,8'h00,
8'h00,8'h07,8'hE0,8'h00,8'hFF,8'hE0,8'h00,8'h00,8'h07,8'h07,8'hE0,8'h01,8'hFF,8'hF8,8'h00,8'h00,
8'h0F,8'hFF,8'hFF,8'h03,8'hFB,8'hFE,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'h87,8'hF0,8'hFF,8'hC0,8'h00,
8'h1F,8'hFF,8'hFF,8'h9F,8'hC0,8'h7F,8'hF0,8'h00,8'h1F,8'hFF,8'hE0,8'h3F,8'h80,8'h1F,8'hFE,8'h00,
8'h08,8'h07,8'hE0,8'hFE,8'h00,8'h0F,8'hFF,8'hC0,8'h00,8'h07,8'hE3,8'hF9,8'hC0,8'h03,8'hFF,8'hF8,
8'h00,8'h07,8'hF3,8'hF3,8'hFF,8'hF9,8'hFF,8'hFC,8'h00,8'h0F,8'hF9,8'hC7,8'hFF,8'hFC,8'hFF,8'hF8,
8'h00,8'h0F,8'hFC,8'h0F,8'hFF,8'hF8,8'h3F,8'hF0,8'h00,8'h1F,8'hFE,8'h0E,8'h0C,8'h00,8'h1F,8'hE0,
8'h00,8'h3F,8'hFF,8'h00,8'h1E,8'h00,8'h0F,8'h80,8'h00,8'h7F,8'hFF,8'h80,8'h3F,8'h01,8'h00,8'h00,
8'h00,8'hFF,8'hE7,8'h84,8'h3F,8'h03,8'hC0,8'h00,8'h01,8'hFF,8'hE0,8'h9E,8'h3F,8'h07,8'hC0,8'h00,
8'h03,8'hFF,8'hE0,8'h1E,8'h3F,8'h0F,8'hE0,8'h00,8'h07,8'hF7,8'hE0,8'h3F,8'h1F,8'h0F,8'hE0,8'h00,
8'h1F,8'hE7,8'hE0,8'h3F,8'h1F,8'h0F,8'hC0,8'h00,8'h3F,8'hC7,8'hE0,8'h1F,8'h0F,8'h0F,8'hC0,8'h00,
8'h7F,8'h87,8'hE0,8'h1F,8'h8F,8'h0F,8'h80,8'h00,8'h7F,8'h07,8'hE0,8'h0F,8'h87,8'h0F,8'h80,8'h00,
8'h3E,8'h07,8'hE0,8'h07,8'h83,8'h1F,8'h00,8'h00,8'h08,8'h07,8'hE0,8'h03,8'hC0,8'h1E,8'h00,8'h00,
8'h00,8'h07,8'hE0,8'h01,8'hC0,8'h1E,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h18,8'hC0,8'h3C,8'h00,8'h00,
8'h00,8'h07,8'hE0,8'h7E,8'h00,8'h38,8'h00,8'h00,8'h00,8'h07,8'hE0,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,
8'h00,8'h07,8'hE1,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h07,8'hE3,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,
8'h00,8'h07,8'hE3,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'h00,8'h07,8'hE3,8'hC0,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "检"
    char[20]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h07,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h60,8'h07,8'hE0,8'h00,8'h00,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,
8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h01,8'h00,8'h0F,8'hE0,8'h00,8'h00,8'h00,
8'h00,8'h20,8'h00,8'h0F,8'hE0,8'h00,8'h00,8'h00,8'h00,8'hF8,8'h00,8'h0F,8'hE0,8'h00,8'h1E,8'h00,
8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,
8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h03,8'hF0,8'h00,8'h0F,8'h00,8'h00,8'h1F,8'h00,
8'h03,8'hE0,8'h00,8'h1F,8'h80,8'h00,8'h0F,8'h00,8'h03,8'hE0,8'h00,8'hFF,8'h03,8'hC0,8'h0F,8'h00,
8'h03,8'hC0,8'h1F,8'hFC,8'h0F,8'hE0,8'h0F,8'h00,8'h01,8'hC0,8'h3F,8'hF0,8'h3F,8'hE0,8'h07,8'h00,
8'h01,8'hC0,8'h7F,8'hF0,8'hFF,8'hC0,8'h07,8'h00,8'h01,8'hC0,8'h7F,8'hFF,8'hFC,8'h00,8'h07,8'h00,
8'h01,8'hC0,8'h20,8'hFF,8'hE0,8'h00,8'h07,8'h00,8'h00,8'hC0,8'h00,8'h3F,8'h01,8'hE0,8'h06,8'h00,
8'h00,8'h00,8'h00,8'hFC,8'h01,8'hF8,8'h06,8'h00,8'h00,8'h00,8'h0F,8'hF0,8'h01,8'hFC,8'h00,8'h00,
8'h00,8'h03,8'hFF,8'hF0,8'h0F,8'hFE,8'h00,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,8'h00,
8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'h1F,8'h00,8'h00,8'h00,8'h03,8'h80,8'h07,8'hE0,8'h0F,8'h80,8'h00,
8'h00,8'h00,8'h0E,8'h03,8'hE0,8'h03,8'h80,8'h00,8'h00,8'h00,8'h1F,8'h03,8'hE1,8'hF1,8'h80,8'h00,
8'h00,8'h00,8'h3F,8'h83,8'hE3,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h7F,8'h03,8'hE3,8'hFC,8'h00,8'h00,
8'h00,8'h01,8'hFE,8'h03,8'hE1,8'hFF,8'h00,8'h00,8'h00,8'h07,8'hF8,8'h03,8'hE0,8'hFF,8'hC0,8'h00,
8'h00,8'h3F,8'hE0,8'h07,8'hE0,8'h1F,8'hF8,8'h00,8'h00,8'hFF,8'h81,8'h87,8'hE0,8'h07,8'hFE,8'h00,
8'h03,8'hFE,8'h01,8'hFF,8'hE0,8'h00,8'h7F,8'h80,8'h00,8'h00,8'h00,8'hFF,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h7F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F,8'h80,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "索"
    char[21]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h1E,8'h00,8'h10,8'h00,8'h07,8'h80,8'h00,8'h00,8'h3F,8'h00,8'h7C,8'h00,8'h1F,8'hC0,8'h00,
8'h00,8'h3F,8'h80,8'h7F,8'h3F,8'hFF,8'hC0,8'h00,8'h00,8'h3F,8'hE0,8'h7F,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h1F,8'hF0,8'h7F,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'h03,8'hF8,8'h7E,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h7C,8'h00,8'h1C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'hE1,8'hFE,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h7D,8'hFF,8'hFE,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3D,8'hFF,8'hBE,8'h00,8'h00,
8'h00,8'hE0,8'h60,8'h3D,8'hE0,8'h1E,8'h00,8'h00,8'h01,8'hFF,8'hF0,8'h3C,8'h00,8'h3E,8'h00,8'h00,
8'h01,8'hFF,8'hF0,8'h3C,8'h00,8'h1C,8'h00,8'h00,8'h01,8'hFF,8'hF0,8'h38,8'h38,8'h3C,8'h00,8'h00,
8'h01,8'h81,8'hE0,8'h38,8'h7C,8'h38,8'h00,8'h00,8'h00,8'h01,8'hC0,8'h38,8'h3F,8'h78,8'h00,8'h00,
8'h00,8'h01,8'h80,8'h78,8'h3F,8'hF0,8'h00,8'h00,8'h00,8'h03,8'h80,8'h78,8'h1F,8'hF0,8'h00,8'h00,
8'h00,8'h03,8'h80,8'hF0,8'h07,8'hF0,8'h00,8'h00,8'h00,8'h03,8'h80,8'hF0,8'h07,8'hF8,8'h00,8'h00,
8'h00,8'h03,8'hC1,8'hE0,8'h1F,8'hFC,8'h00,8'h00,8'h00,8'h01,8'hC7,8'hC0,8'hFF,8'hFE,8'h00,8'h00,
8'h00,8'h01,8'hCF,8'h9F,8'hFE,8'h3F,8'h00,8'h00,8'h00,8'h01,8'hC7,8'h3F,8'hF8,8'h1F,8'h80,8'h00,
8'h00,8'h03,8'h80,8'h1F,8'hE0,8'h07,8'hC0,8'h00,8'h01,8'hFF,8'h80,8'h00,8'h00,8'h03,8'hE0,8'h00,
8'h0F,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'hF8,8'h00,8'h1F,8'hFF,8'hFC,8'h00,8'h00,8'h00,8'h78,8'h00,
8'h3F,8'hFF,8'hFF,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h3F,8'hE3,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h02,
8'h3E,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h38,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,
8'h00,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'hF0,
8'h00,8'h00,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hC0,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hFF,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "返"
    char[22]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h10,8'h00,
8'h00,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'h7C,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,
8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,
8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,8'h00,8'hFE,8'h00,8'h00,8'h00,8'h00,8'hFE,8'h00,
8'h00,8'h7E,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,
8'h00,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h7C,8'h0F,8'hE0,8'h03,8'hC0,8'h7E,8'h00,
8'h00,8'h7C,8'h0F,8'hFF,8'hFF,8'hE0,8'h7E,8'h00,8'h00,8'h7C,8'h1F,8'hFF,8'hFF,8'hE0,8'h7C,8'h00,
8'h00,8'h7C,8'h0F,8'hFF,8'hFF,8'hE0,8'h7C,8'h00,8'h00,8'h7C,8'h0F,8'h80,8'h07,8'hE0,8'h7C,8'h00,
8'h00,8'h7C,8'h0F,8'h80,8'h07,8'hE0,8'h7C,8'h00,8'h00,8'h7C,8'h0F,8'h80,8'h07,8'hE0,8'h7C,8'h00,
8'h00,8'h7C,8'h0F,8'h80,8'h07,8'hE0,8'h7C,8'h00,8'h00,8'h7C,8'h0F,8'h80,8'h07,8'hE0,8'h7C,8'h00,
8'h00,8'h7C,8'h0F,8'h80,8'h07,8'hE0,8'h7C,8'h00,8'h00,8'h7C,8'h0F,8'hFF,8'hEF,8'hE0,8'h7C,8'h00,
8'h00,8'h7C,8'h07,8'hFF,8'hFF,8'hE0,8'h7C,8'h00,8'h00,8'h7C,8'h07,8'hFF,8'hFF,8'hC0,8'h7C,8'h00,
8'h00,8'h7C,8'h07,8'hFF,8'hFF,8'hC0,8'hFC,8'h00,8'h00,8'h7C,8'h07,8'h80,8'h07,8'hC0,8'hFC,8'h00,
8'h00,8'h7E,8'h00,8'h00,8'h01,8'h00,8'hFC,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,8'h00,8'hFC,8'h00,
8'h00,8'h7E,8'h00,8'h00,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,8'h01,8'hFC,8'h00,
8'h00,8'h7F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,
8'h00,8'h7F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,
8'h00,8'h7F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h18,8'h00,8'h00,8'h00,8'h00,8'hF8,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "回"
    char[23]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h07,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hE0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,
8'h00,8'h7F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'hFF,8'hF8,8'h0F,8'hFF,8'hFF,8'hFF,8'h00,
8'h00,8'hFC,8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h00,8'hE1,8'h80,8'h3E,8'h00,8'h0E,8'h00,8'h00,
8'h00,8'h07,8'hC1,8'hFC,8'h30,8'h1E,8'h00,8'h00,8'h00,8'h07,8'hE1,8'hF0,8'h7C,8'h3E,8'h00,8'h00,
8'h00,8'h07,8'hF3,8'hF8,8'hF8,8'h7C,8'h00,8'h00,8'h00,8'h03,8'hFB,8'hFF,8'hF8,8'hF8,8'h00,8'h00,
8'h00,8'h00,8'h71,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h00,8'hF0,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h1E,8'h38,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h1C,8'h3C,8'h3C,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'hFD,8'hFC,8'h1E,8'h7E,8'h00,8'h00,8'h00,8'h0F,8'hF9,8'hFF,8'hFF,8'h3F,8'h80,8'h00,
8'h00,8'h1F,8'hF1,8'hFF,8'hE3,8'h0F,8'hE0,8'h00,8'h00,8'h1F,8'hC0,8'h1F,8'hC1,8'h01,8'hE0,8'h00,
8'h00,8'h0F,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,
8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,
8'h3F,8'hFF,8'hF0,8'h0F,8'hFF,8'hFF,8'hFF,8'hF0,8'h3F,8'hC0,8'h00,8'h0F,8'hC0,8'h0F,8'hFF,8'hE0,
8'h3C,8'h00,8'h00,8'h0F,8'hC0,8'h01,8'hFF,8'h80,8'h10,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h3E,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "律"
    char[24]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F,8'hFF,8'hF8,8'h00,
8'h3F,8'hFF,8'hFF,8'h00,8'h07,8'hE0,8'h1F,8'hC0,8'h03,8'hC0,8'h07,8'hE0,8'h03,8'hC0,8'h03,8'hF0,
8'h03,8'hC0,8'h01,8'hF0,8'h03,8'hC0,8'h01,8'hF8,8'h03,8'hC0,8'h00,8'hF8,8'h03,8'hC0,8'h00,8'hF8,
8'h03,8'hC0,8'h00,8'hF8,8'h03,8'hC0,8'h00,8'hF8,8'h03,8'hC0,8'h00,8'hF8,8'h03,8'hC0,8'h00,8'hF8,
8'h03,8'hC0,8'h00,8'hF8,8'h03,8'hC0,8'h01,8'hF0,8'h03,8'hC0,8'h01,8'hF0,8'h03,8'hC0,8'h03,8'hE0,
8'h03,8'hC0,8'h07,8'hC0,8'h03,8'hC0,8'h1F,8'h80,8'h03,8'hFF,8'hFF,8'h00,8'h03,8'hFF,8'hF8,8'h00,
8'h03,8'hC0,8'hF0,8'h00,8'h03,8'hC0,8'hF8,8'h00,8'h03,8'hC0,8'h78,8'h00,8'h03,8'hC0,8'h7C,8'h00,
8'h03,8'hC0,8'h3C,8'h00,8'h03,8'hC0,8'h3C,8'h00,8'h03,8'hC0,8'h3E,8'h00,8'h03,8'hC0,8'h1E,8'h00,
8'h03,8'hC0,8'h1F,8'h00,8'h03,8'hC0,8'h0F,8'h00,8'h03,8'hC0,8'h0F,8'h80,8'h03,8'hC0,8'h07,8'h80,
8'h03,8'hC0,8'h07,8'h80,8'h03,8'hC0,8'h07,8'hC0,8'h03,8'hC0,8'h03,8'hC0,8'h03,8'hC0,8'h03,8'hE0,
8'h03,8'hC0,8'h01,8'hE0,8'h03,8'hC0,8'h01,8'hE0,8'h03,8'hC0,8'h00,8'hF0,8'h07,8'hE0,8'h00,8'hF8,
8'h3F,8'hFC,8'h00,8'hFF,8'h3F,8'hFC,8'h00,8'h7F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "R"
    char[25]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3C,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h7E,8'h01,8'hC0,8'h00,8'h18,8'h00,8'h00,8'h00,8'h3F,8'h03,8'hFE,8'h07,8'hFC,8'h00,
8'h00,8'h00,8'h1F,8'h87,8'hFF,8'hFF,8'hFE,8'h00,8'h00,8'h00,8'h07,8'hC7,8'hFF,8'hFF,8'hFE,8'h00,
8'h00,8'h1C,8'h00,8'h07,8'hC0,8'h07,8'hFE,8'h00,8'h00,8'h1E,8'h00,8'h06,8'h00,8'h00,8'hFE,8'h00,
8'h00,8'h1E,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'hFE,8'h00,
8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'hFE,8'h00,8'h00,8'h1F,8'h03,8'h00,8'h00,8'h00,8'hFC,8'h00,
8'h00,8'h0F,8'h07,8'hFF,8'hFF,8'hE0,8'hFC,8'h00,8'h00,8'h0F,8'h07,8'hFF,8'hFF,8'hE0,8'hFC,8'h00,
8'h00,8'h0F,8'h07,8'hFF,8'hFF,8'hE0,8'hFC,8'h00,8'h00,8'h0F,8'h07,8'hC0,8'h07,8'hE0,8'hFC,8'h00,
8'h00,8'h0F,8'h07,8'hC0,8'h03,8'hE0,8'hFC,8'h00,8'h00,8'h0F,8'h07,8'h80,8'h03,8'hE0,8'hFC,8'h00,
8'h00,8'h1F,8'h07,8'h80,8'h03,8'hE0,8'hFC,8'h00,8'h00,8'h1F,8'h07,8'hC0,8'h07,8'hE0,8'hFC,8'h00,
8'h00,8'h1F,8'h07,8'hFF,8'hFF,8'hE0,8'hFC,8'h00,8'h00,8'h1F,8'h03,8'hFF,8'hFF,8'hE0,8'hFC,8'h00,
8'h00,8'h1F,8'h03,8'hFF,8'hFF,8'hE0,8'hFC,8'h00,8'h00,8'h3F,8'h03,8'hC0,8'h03,8'hE0,8'hFC,8'h00,
8'h00,8'h3E,8'h03,8'hC0,8'h03,8'hE0,8'hFC,8'h00,8'h00,8'h7E,8'h03,8'hC0,8'h03,8'hE0,8'hFC,8'h00,
8'h00,8'h7E,8'h03,8'hC0,8'h03,8'hE0,8'hFE,8'h00,8'h00,8'hFE,8'h03,8'hC0,8'h03,8'hE0,8'hFE,8'h00,
8'h01,8'hFC,8'h03,8'hFF,8'hFF,8'hE0,8'hFE,8'h00,8'h03,8'hFC,8'h03,8'hFF,8'hFF,8'hE0,8'hFE,8'h00,
8'h07,8'hFC,8'h03,8'hFF,8'hFF,8'hE0,8'hFE,8'h00,8'h3F,8'hF8,8'h01,8'hC0,8'h01,8'h80,8'hFE,8'h00,
8'h3F,8'hF0,8'h00,8'h00,8'h00,8'h00,8'hFE,8'h00,8'h3F,8'hF0,8'h00,8'h00,8'h00,8'h00,8'hFF,8'h00,
8'h3F,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h7F,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "间"
    char[26]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0E,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hE0,8'h1F,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h01,8'hF0,8'h1F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h01,8'hF0,8'h1F,8'h80,8'hF0,8'h0E,8'h00,
8'h00,8'h01,8'hF0,8'h1F,8'h81,8'hFF,8'hFF,8'h80,8'h00,8'h01,8'hF0,8'h1F,8'h81,8'hFF,8'hFF,8'h80,
8'h00,8'hFF,8'hFF,8'hFF,8'hF1,8'hFF,8'hFF,8'h80,8'h01,8'hFF,8'hFF,8'hFF,8'hF9,8'hFF,8'hFF,8'h80,
8'h01,8'hFF,8'hFF,8'hFF,8'hF1,8'hF0,8'h1F,8'h80,8'h01,8'hE1,8'hF0,8'h0F,8'h01,8'hE0,8'h0F,8'h80,
8'h00,8'h01,8'hF0,8'h0F,8'h01,8'hE0,8'h0F,8'h80,8'h00,8'h01,8'hF9,8'hFF,8'h01,8'hE0,8'h0F,8'h80,
8'h00,8'h01,8'hFF,8'hFF,8'h01,8'hF0,8'h1F,8'h80,8'h00,8'h01,8'hFF,8'hFF,8'h01,8'hFF,8'hFF,8'h80,
8'h00,8'h01,8'hF0,8'h3F,8'h01,8'hFF,8'hFF,8'h80,8'h00,8'h01,8'hF0,8'h0F,8'h01,8'hFF,8'hFF,8'h80,
8'h00,8'h01,8'hF8,8'h0F,8'h01,8'hFF,8'h3F,8'h80,8'h00,8'h01,8'hFF,8'hFF,8'h01,8'hF0,8'h1F,8'h80,
8'h00,8'h01,8'hFF,8'hFF,8'h01,8'hE0,8'h0F,8'h80,8'h00,8'h01,8'hFF,8'hFF,8'h01,8'hE0,8'h0F,8'h80,
8'h00,8'h01,8'hF0,8'h0F,8'h01,8'hE0,8'h0F,8'h80,8'h00,8'h01,8'hF0,8'h0F,8'h01,8'hF0,8'h1F,8'h80,
8'h00,8'h01,8'hF8,8'h0F,8'h01,8'hFF,8'hFF,8'h80,8'h0F,8'hFF,8'hFF,8'hFF,8'hFD,8'hFF,8'hFF,8'h80,
8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h1F,8'h80,
8'h3F,8'hFF,8'hFF,8'hFF,8'hE3,8'hC0,8'h1F,8'h80,8'h3F,8'h80,8'h00,8'h00,8'h07,8'hC0,8'h1F,8'h80,
8'h38,8'h00,8'h70,8'h1C,8'h07,8'hC0,8'h1F,8'h80,8'h00,8'h00,8'hF8,8'h3E,8'h0F,8'h80,8'h1F,8'h80,
8'h00,8'h01,8'hF8,8'h3F,8'h1F,8'h80,8'h1F,8'h80,8'h00,8'h03,8'hF8,8'h3F,8'hBF,8'h80,8'h1F,8'h80,
8'h00,8'h03,8'hF0,8'h0F,8'hFF,8'h00,8'h1F,8'h80,8'h00,8'h07,8'hE0,8'h00,8'hFE,8'h00,8'h1F,8'h80,
8'h00,8'h0F,8'h80,8'h03,8'hFE,8'h00,8'h1F,8'hC0,8'h00,8'h1F,8'h00,8'h1F,8'hFC,8'h00,8'h1F,8'hC0,
8'h00,8'h3E,8'h00,8'h3F,8'hF8,8'h00,8'h1F,8'hC0,8'h00,8'hF8,8'h00,8'h3F,8'hF0,8'h00,8'h1F,8'hC0,
8'h00,8'hF0,8'h00,8'h0F,8'h80,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "期"
    char[27]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h7F,8'hF8,8'h0F,8'hFF,8'h7F,8'hF8,8'h0F,8'hFF,8'h0F,8'hC0,8'h01,8'hF8,8'h07,8'h80,8'h00,8'hF0,
8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,
8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,
8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,
8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,
8'h07,8'hFF,8'hFF,8'hF0,8'h07,8'hFF,8'hFF,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,
8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,
8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,
8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,
8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF0,
8'h0F,8'hC0,8'h01,8'hF8,8'h7F,8'hF8,8'h0F,8'hFF,8'h7F,8'hF8,8'h0F,8'hFF,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "H"
    char[28]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h7F,8'hF0,8'h03,8'hFE,8'h7F,8'hF0,8'h03,8'hFE,8'h0F,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'h60,
8'h07,8'h80,8'h00,8'h60,8'h07,8'h80,8'h00,8'h60,8'h07,8'hC0,8'h00,8'hC0,8'h03,8'hC0,8'h00,8'hC0,
8'h03,8'hC0,8'h00,8'hC0,8'h03,8'hC0,8'h00,8'hC0,8'h03,8'hE0,8'h01,8'h80,8'h01,8'hE0,8'h01,8'h80,
8'h01,8'hE0,8'h01,8'h80,8'h01,8'hE0,8'h01,8'h80,8'h01,8'hF0,8'h03,8'h00,8'h00,8'hF0,8'h03,8'h00,
8'h00,8'hF0,8'h03,8'h00,8'h00,8'hF0,8'h07,8'h00,8'h00,8'h78,8'h06,8'h00,8'h00,8'h78,8'h06,8'h00,
8'h00,8'h78,8'h06,8'h00,8'h00,8'h78,8'h0E,8'h00,8'h00,8'h3C,8'h0C,8'h00,8'h00,8'h3C,8'h0C,8'h00,
8'h00,8'h3C,8'h0C,8'h00,8'h00,8'h3E,8'h18,8'h00,8'h00,8'h1E,8'h18,8'h00,8'h00,8'h1E,8'h18,8'h00,
8'h00,8'h1E,8'h18,8'h00,8'h00,8'h1F,8'h30,8'h00,8'h00,8'h0F,8'h30,8'h00,8'h00,8'h0F,8'h30,8'h00,
8'h00,8'h0F,8'h30,8'h00,8'h00,8'h0F,8'hE0,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h00,8'h07,8'hE0,8'h00,
8'h00,8'h07,8'hE0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h01,8'h80,8'h00,8'h00,8'h01,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "V"
    char[29]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h78,8'h00,8'h3C,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFC,8'h00,8'h3F,8'h00,8'h00,8'h00,
8'h00,8'h00,8'hFC,8'h00,8'h3F,8'h00,8'h60,8'h00,8'h00,8'h00,8'hFE,8'h00,8'h3F,8'h00,8'hF0,8'h00,
8'h00,8'h00,8'hFE,8'h00,8'h3F,8'h01,8'hF0,8'h00,8'h00,8'h00,8'hFE,8'h00,8'h3F,8'h03,8'hF0,8'h00,
8'h07,8'h80,8'hFE,8'h00,8'h3F,8'h07,8'hE0,8'h00,8'h0F,8'hC0,8'hFE,8'h00,8'h3F,8'h0F,8'h80,8'h00,
8'h0F,8'hE0,8'hFE,8'h00,8'h3F,8'h0E,8'h00,8'h00,8'h07,8'hF0,8'h7E,8'h00,8'h3F,8'h00,8'h00,8'h00,
8'h03,8'hF0,8'h7E,8'h00,8'h3F,8'h00,8'h00,8'h00,8'h01,8'hF8,8'h7E,8'h20,8'h3F,8'h00,8'h00,8'h00,
8'h00,8'hFC,8'h7E,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h3E,8'h7E,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,
8'h00,8'h0F,8'h7F,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h7F,8'h80,8'h3F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h3F,8'hC0,8'h00,8'h00,
8'h00,8'h01,8'hFE,8'h00,8'h7F,8'hE0,8'h00,8'h00,8'h00,8'h07,8'hFE,8'h00,8'h7F,8'hF0,8'h00,8'h00,
8'h00,8'h1F,8'hFE,8'h00,8'hFD,8'hF8,8'h00,8'h00,8'h00,8'hFF,8'h7E,8'h00,8'hF8,8'hFC,8'h00,8'h00,
8'h0F,8'hFE,8'h7E,8'h01,8'hF8,8'h7F,8'h00,8'h00,8'h1F,8'hFC,8'h7E,8'h01,8'hF8,8'h3F,8'h80,8'h00,
8'h3F,8'hF8,8'h7E,8'h03,8'hF0,8'h1F,8'hC0,8'h00,8'h3F,8'hE0,8'h7E,8'h03,8'hF0,8'h0F,8'hF0,8'h00,
8'h3F,8'hC0,8'h7E,8'h07,8'hE0,8'h07,8'hF8,8'h00,8'h3F,8'h00,8'h7E,8'h0F,8'hE0,8'h03,8'hFE,8'h00,
8'h1E,8'h00,8'h7E,8'h1F,8'hC0,8'h03,8'hFF,8'h00,8'h00,8'h00,8'h7E,8'h3F,8'h80,8'h01,8'hFF,8'hC0,
8'h00,8'h00,8'h7E,8'h7F,8'h00,8'h00,8'hFF,8'hF0,8'h00,8'h00,8'h7F,8'hFE,8'h00,8'h00,8'h7F,8'hFC,
8'h00,8'h00,8'hFF,8'hFC,8'h00,8'h00,8'h7F,8'hFC,8'h00,8'h00,8'hFF,8'hF0,8'h00,8'h00,8'h3F,8'hFC,
8'h00,8'h00,8'hFE,8'h00,8'h00,8'h00,8'h1F,8'hF8,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h1F,8'hF0,
8'h00,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h70,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "状"
    char[30]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h1F,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hE0,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h01,8'h80,8'h3E,8'h3E,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h7C,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'hFC,8'h0F,8'hC0,8'h00,8'h00,
8'h00,8'h00,8'h03,8'hFA,8'h07,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hE7,8'h03,8'hF8,8'h00,8'h00,
8'h00,8'h00,8'hFF,8'hC7,8'h81,8'hFE,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'h87,8'hE0,8'h7F,8'h00,8'h00,
8'h00,8'h3F,8'hFE,8'h07,8'hF0,8'h3F,8'hC0,8'h00,8'h00,8'h0F,8'hF8,8'h00,8'h20,8'h0F,8'hF0,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h18,8'h78,8'h00,
8'h00,8'h00,8'h1C,8'h00,8'h78,8'h3C,8'h00,8'h00,8'h00,8'h04,8'h1F,8'h00,8'h7C,8'h7E,8'h00,8'h00,
8'h00,8'h04,8'h3F,8'h80,8'hF8,8'h7E,8'h00,8'h00,8'h00,8'h0C,8'h3F,8'hE0,8'hF0,8'hFC,8'h00,8'h00,
8'h00,8'h1C,8'h3F,8'hF0,8'hE1,8'hFC,8'h00,8'h00,8'h00,8'h3C,8'h38,8'hFD,8'hC1,8'hF8,8'h00,8'h00,
8'h00,8'h7C,8'h30,8'h7F,8'h83,8'hF0,8'h00,8'h00,8'h00,8'hF8,8'h00,8'h3F,8'hC7,8'hC0,8'h00,8'h00,
8'h01,8'hF8,8'h00,8'h0F,8'hFF,8'h00,8'h00,8'h00,8'h03,8'hF8,8'h00,8'h07,8'hFC,8'h00,8'h00,8'h02,
8'h07,8'hF8,8'h00,8'h01,8'hFF,8'hF8,8'h00,8'hFC,8'h0F,8'hF0,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hF8,
8'h0F,8'hF0,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'hF8,8'h0F,8'hE0,8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hF0,
8'h0F,8'hC0,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hE0,8'h0F,8'hC0,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hC0,
8'h00,8'h00,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F,8'hFF,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hFE,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'hF0,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "态"
    char[31]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,
8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,
8'h00,8'h1F,8'hF0,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h1F,8'h00,8'h03,8'hF8,8'h00,8'h00,8'h00,
8'h00,8'h1C,8'h00,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hF8,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hF8,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hF8,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h78,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7C,8'h03,8'hFF,8'hF8,8'h00,8'h00,
8'h00,8'h00,8'h7E,8'h03,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h03,8'hFF,8'hFF,8'h80,8'h00,
8'h00,8'h00,8'h7E,8'h03,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h03,8'hFF,8'hFE,8'h00,8'h00,
8'h00,8'h00,8'h3E,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h03,8'hF8,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h3E,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h03,8'hF8,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h3E,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h03,8'hF8,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h3E,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h03,8'hF8,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h3E,8'h03,8'hF8,8'h00,8'h00,8'h00,8'h02,8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hE0,8'h04,
8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,
8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h3F,8'hFF,8'hFF,8'hC0,8'h7F,8'hFF,8'hFF,8'hF8,
8'h3F,8'hFE,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hF0,8'h3F,8'hC0,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hF0,
8'h1C,8'h00,8'h00,8'h00,8'h00,8'h01,8'hFF,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F,8'hC0,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "正"
    char[32]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h08,8'h0F,8'hC0,8'h38,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h0F,8'hE0,8'h7C,8'h00,8'h00,
8'h00,8'h00,8'h7E,8'h0F,8'hC0,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h7F,8'h0F,8'hC0,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'h7F,8'h0F,8'hC0,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h3F,8'h0F,8'hC1,8'hF0,8'h00,8'h00,
8'h00,8'h00,8'h0F,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'hF0,8'h00,8'h0F,8'hC0,8'h00,8'h3F,8'h80,
8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,
8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h03,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hE0,
8'h03,8'hF0,8'h0E,8'h00,8'h00,8'hC0,8'h03,8'hE0,8'h03,8'hE0,8'h1F,8'hFF,8'hFF,8'hE0,8'h03,8'hE0,
8'h03,8'hE0,8'h1F,8'hFF,8'hFF,8'hF0,8'h01,8'hE0,8'h03,8'hC0,8'h1F,8'hFF,8'hFF,8'hF0,8'h01,8'hE0,
8'h03,8'hC0,8'h1F,8'h00,8'h01,8'hF0,8'h01,8'hE0,8'h03,8'hC0,8'h1F,8'h00,8'h01,8'hF0,8'h01,8'hC0,
8'h01,8'hC0,8'h1F,8'hFF,8'hFF,8'hF0,8'h01,8'hC0,8'h01,8'h80,8'h1F,8'hFF,8'hFF,8'hE0,8'h00,8'hC0,
8'h00,8'h80,8'h0F,8'hFF,8'hFF,8'hE0,8'h00,8'h80,8'h00,8'h00,8'h04,8'h0F,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h40,8'h0F,8'hC0,8'h07,8'h80,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'hF0,8'h0F,8'hC0,8'h1F,8'hC0,8'h00,
8'h00,8'h00,8'hF0,8'h0F,8'hC0,8'h1F,8'hC0,8'h00,8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h03,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h07,8'hE0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h0F,8'hE0,8'h0F,8'hC0,8'h1F,8'hC0,8'h00,
8'h00,8'h0F,8'hC0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h0F,8'h00,8'h0F,8'hC0,8'h0F,8'h80,8'h00,
8'h00,8'h00,8'h00,8'h07,8'h80,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "常"
    char[33]  <= {
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h08,8'h0F,8'hC0,8'h38,8'h00,8'h00,8'h00,8'h00,8'h3E,8'h0F,8'hE0,8'h7C,8'h00,8'h00,
8'h00,8'h00,8'h7E,8'h0F,8'hC0,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h7F,8'h0F,8'hC0,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'h7F,8'h0F,8'hC0,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h3F,8'h0F,8'hC1,8'hF0,8'h00,8'h00,
8'h00,8'h00,8'h0F,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'hF0,8'h00,8'h0F,8'hC0,8'h00,8'h3F,8'h80,
8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,
8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h03,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hE0,
8'h03,8'hF0,8'h0E,8'h00,8'h00,8'hC0,8'h03,8'hE0,8'h03,8'hE0,8'h1F,8'hFF,8'hFF,8'hE0,8'h03,8'hE0,
8'h03,8'hE0,8'h1F,8'hFF,8'hFF,8'hF0,8'h01,8'hE0,8'h03,8'hC0,8'h1F,8'hFF,8'hFF,8'hF0,8'h01,8'hE0,
8'h03,8'hC0,8'h1F,8'h00,8'h01,8'hF0,8'h01,8'hE0,8'h03,8'hC0,8'h1F,8'h00,8'h01,8'hF0,8'h01,8'hC0,
8'h01,8'hC0,8'h1F,8'hFF,8'hFF,8'hF0,8'h01,8'hC0,8'h01,8'h80,8'h1F,8'hFF,8'hFF,8'hE0,8'h00,8'hC0,
8'h00,8'h80,8'h0F,8'hFF,8'hFF,8'hE0,8'h00,8'h80,8'h00,8'h00,8'h04,8'h0F,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h40,8'h0F,8'hC0,8'h07,8'h80,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'hF0,8'h0F,8'hC0,8'h1F,8'hC0,8'h00,
8'h00,8'h00,8'hF0,8'h0F,8'hC0,8'h1F,8'hC0,8'h00,8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h03,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h07,8'hE0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h0F,8'hE0,8'h0F,8'hC0,8'h1F,8'hC0,8'h00,
8'h00,8'h0F,8'hC0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h0F,8'h00,8'h0F,8'hC0,8'h0F,8'h80,8'h00,
8'h00,8'h00,8'h00,8'h07,8'h80,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "轻"
    char[34]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hE0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h03,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hF0,8'h00,8'h00,8'h00,
8'h00,8'h03,8'h80,8'h07,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h07,8'hF0,8'h07,8'hFF,8'hC0,8'h00,8'h00,
8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,
8'h00,8'h07,8'hC0,8'h7C,8'h01,8'hFF,8'hF0,8'h00,8'h00,8'h07,8'h80,8'h3C,8'h01,8'hE0,8'h00,8'h00,
8'h00,8'h07,8'h80,8'h3C,8'h01,8'hE0,8'h00,8'h00,8'h00,8'h07,8'h80,8'h3C,8'h01,8'hE0,8'h00,8'h00,
8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,
8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h07,8'hC0,8'h3C,8'h01,8'hE0,8'h00,8'h00,
8'h00,8'h07,8'h80,8'h3C,8'h01,8'hE0,8'h00,8'h00,8'h00,8'h07,8'h80,8'h3C,8'h03,8'hE0,8'h00,8'h00,
8'h00,8'h07,8'h80,8'h3F,8'hFF,8'hE0,8'h00,8'h00,8'h00,8'h07,8'h80,8'h3F,8'hFF,8'hE0,8'h00,8'h00,
8'h00,8'h07,8'h80,8'h3E,8'h07,8'hE0,8'h00,8'h00,8'h00,8'h07,8'h80,8'h00,8'h00,8'hC0,8'h00,8'h00,
8'h00,8'h0F,8'h80,8'h21,8'hFE,8'h30,8'h00,8'h00,8'h00,8'h0F,8'h80,8'hFF,8'hFF,8'hF8,8'h00,8'h00,
8'h00,8'h1F,8'h80,8'hFF,8'hFF,8'hF8,8'h00,8'h00,8'h00,8'h1F,8'h00,8'hFE,8'h01,8'hF8,8'h00,8'h00,
8'h00,8'h3F,8'h00,8'hFF,8'h01,8'hF0,8'h00,8'h00,8'h00,8'h3F,8'h00,8'h1F,8'hE3,8'hE0,8'h00,8'h00,
8'h00,8'h7E,8'h00,8'h07,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'hFE,8'h00,8'h01,8'hFF,8'hC0,8'h00,8'h00,
8'h01,8'hFE,8'h00,8'h00,8'h7F,8'h80,8'h00,8'h00,8'h03,8'hFC,8'h00,8'h00,8'h3F,8'hF0,8'h00,8'h00,
8'h0F,8'hF8,8'h00,8'h00,8'h7F,8'hFF,8'h00,8'h00,8'h1F,8'hF8,8'h00,8'h01,8'hFF,8'hFF,8'hF0,8'h00,
8'h3F,8'hF0,8'h00,8'h0F,8'hF0,8'hFF,8'hFF,8'hE2,8'h1F,8'hE0,8'h00,8'hFF,8'hE0,8'h3F,8'hFF,8'hFC,
8'h1F,8'hC3,8'hFF,8'hFF,8'h80,8'h0F,8'hFF,8'hFC,8'h00,8'h01,8'hFF,8'hFE,8'h00,8'h03,8'hFF,8'hF8,
8'h00,8'h01,8'hFF,8'hF0,8'h00,8'h00,8'hFF,8'hF0,8'h00,8'h00,8'hFF,8'h80,8'h00,8'h00,8'h7F,8'hF0,
8'h00,8'h00,8'h30,8'h00,8'h00,8'h00,8'h1F,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "度"
    char[35]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hE0,8'h00,
8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,
8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h06,8'h00,8'h3C,8'h3E,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h18,8'h3C,8'h3E,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h3C,8'h3C,8'h3E,8'h1F,8'h00,8'h00,
8'h00,8'h00,8'h3E,8'h3C,8'h3E,8'h3F,8'h00,8'h00,8'h00,8'h00,8'h3F,8'h3C,8'h3E,8'h3E,8'h00,8'h00,
8'h00,8'h00,8'h3F,8'h3C,8'h3E,8'h7E,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hBC,8'h3E,8'hF8,8'h00,8'h00,
8'h00,8'h00,8'h01,8'h3C,8'h3E,8'h40,8'h00,8'h00,8'h00,8'h07,8'h80,8'h3E,8'h3E,8'h00,8'h00,8'h00,
8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,
8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,8'h3F,8'hFF,8'hC0,8'h1F,8'hFF,8'hFF,8'hF0,
8'h00,8'h1F,8'hE0,8'h00,8'h00,8'h0F,8'hFF,8'hE0,8'h00,8'h1F,8'hC0,8'h00,8'h00,8'h00,8'hFF,8'hC0,
8'h00,8'h1F,8'h80,8'h00,8'h00,8'h00,8'h1F,8'h80,8'h00,8'h1F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h1F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h3F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'hFE,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'hFE,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h07,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h3F,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h03,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "严"
    char[36]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0C,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h7F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hFF,8'h80,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hF0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h07,8'hF0,8'h00,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFE,
8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,
8'h1F,8'hFE,8'h00,8'h03,8'hF0,8'h3F,8'hFF,8'hF8,8'h1F,8'hC0,8'h20,8'h03,8'hF0,8'h00,8'h7F,8'hF8,
8'h1C,8'h01,8'hF8,8'h07,8'hF0,8'h0F,8'h07,8'hF0,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h03,8'hFC,8'h03,8'hF0,8'h1F,8'hC0,8'h00,
8'h00,8'h01,8'hF8,8'h03,8'hF0,8'h1F,8'hC0,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h01,8'hFC,8'h07,8'hFF,8'hFF,8'h80,8'h00,
8'h00,8'h01,8'hF8,8'h03,8'hF0,8'h1F,8'h80,8'h00,8'h00,8'h00,8'hF8,8'h03,8'hF0,8'h1F,8'h80,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hF0,8'h7F,8'h00,8'h00,8'h00,8'h00,8'hF0,8'h03,8'hF0,8'h06,8'h00,8'h00,
8'h00,8'h00,8'h10,8'h03,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hE0,8'h00,
8'h00,8'h00,8'h60,8'h03,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hF0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h07,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,
8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,
8'h00,8'h3F,8'hE0,8'h00,8'h00,8'h0F,8'hFF,8'hC0,8'h00,8'h1C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "重"
    char[37]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h01,8'hFC,8'h00,8'h00,8'h70,8'h00,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'hF8,8'h00,8'h00,8'h7C,8'h00,8'h00,8'h00,8'h00,8'hF0,8'h00,8'h00,8'h7C,8'h00,8'h00,
8'h00,8'h00,8'hF0,8'h00,8'h00,8'hFC,8'h00,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'h00,
8'h00,8'h01,8'hF8,8'h00,8'h00,8'h78,8'h00,8'h00,8'h00,8'h01,8'hF0,8'h00,8'h00,8'h00,8'h06,8'h00,
8'h00,8'h01,8'hF0,8'h00,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h01,8'hF8,8'h00,8'h00,8'h01,8'hFC,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hE0,8'h00,
8'h00,8'h00,8'h07,8'hE0,8'h01,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h03,8'hC0,8'h00,8'h00,
8'h00,8'h00,8'h07,8'hE0,8'h07,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h07,8'hE0,8'h07,8'hE0,8'h00,8'h00,
8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,
8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,
8'h3F,8'hF0,8'h07,8'hE0,8'h07,8'hE1,8'hFF,8'hF0,8'h3E,8'h00,8'h07,8'hE0,8'h07,8'hE0,8'h0F,8'hE0,
8'h30,8'h00,8'h07,8'hE0,8'h07,8'hE0,8'h03,8'h80,8'h00,8'h00,8'h0F,8'hC0,8'h07,8'hE0,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'hC0,8'h07,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h3F,8'hC0,8'h07,8'hE0,8'h00,8'h00,
8'h00,8'h00,8'h7F,8'h80,8'h07,8'hE0,8'h00,8'h00,8'h00,8'h03,8'hFF,8'h00,8'h07,8'hE0,8'h00,8'h00,
8'h00,8'h7F,8'hFE,8'h00,8'h07,8'hE0,8'h00,8'h00,8'h00,8'h7F,8'hFC,8'h00,8'h07,8'hE0,8'h00,8'h00,
8'h00,8'h3F,8'hF8,8'h00,8'h0F,8'hE0,8'h00,8'h00,8'h00,8'h07,8'hC0,8'h00,8'h07,8'hC0,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "异"
    char[38]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h0F,8'hC0,8'h38,8'h00,8'h00,
8'h00,8'h00,8'h3E,8'h0F,8'hE0,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h0F,8'hC0,8'h7C,8'h00,8'h00,
8'h00,8'h00,8'h7F,8'h0F,8'hC0,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h7F,8'h0F,8'hC0,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'h3F,8'h0F,8'hC1,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h0F,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'hF0,8'h00,8'h0F,8'hC0,8'h00,8'h3F,8'h80,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,
8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,
8'h03,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hE0,8'h03,8'hF0,8'h0E,8'h00,8'h00,8'hC0,8'h03,8'hE0,
8'h03,8'hE0,8'h1F,8'hFF,8'hFF,8'hE0,8'h03,8'hE0,8'h03,8'hE0,8'h1F,8'hFF,8'hFF,8'hF0,8'h01,8'hE0,
8'h03,8'hC0,8'h1F,8'hFF,8'hFF,8'hF0,8'h01,8'hE0,8'h03,8'hC0,8'h1F,8'h00,8'h01,8'hF0,8'h01,8'hE0,
8'h03,8'hC0,8'h1F,8'h00,8'h01,8'hF0,8'h01,8'hC0,8'h01,8'hC0,8'h1F,8'hFF,8'hFF,8'hF0,8'h01,8'hC0,
8'h01,8'h80,8'h1F,8'hFF,8'hFF,8'hE0,8'h00,8'hC0,8'h00,8'h80,8'h0F,8'hFF,8'hFF,8'hE0,8'h00,8'h80,
8'h00,8'h00,8'h04,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h0F,8'hC0,8'h07,8'h80,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h01,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h00,8'h00,8'hF0,8'h0F,8'hC0,8'h1F,8'hC0,8'h00,8'h00,8'h00,8'hF0,8'h0F,8'hC0,8'h1F,8'hC0,8'h00,
8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h01,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h03,8'hF0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,8'h00,8'h07,8'hE0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h0F,8'hE0,8'h0F,8'hC0,8'h1F,8'hC0,8'h00,8'h00,8'h0F,8'hC0,8'h0F,8'hC0,8'h0F,8'hC0,8'h00,
8'h00,8'h0F,8'h00,8'h0F,8'hC0,8'h0F,8'h80,8'h00,8'h00,8'h00,8'h00,8'h07,8'h80,8'h06,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "常"
    char[39]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h7F,8'hFF,8'h80,8'h00,8'h7F,8'hFF,8'hF0,8'h00,8'h0F,8'hC0,8'hFC,8'h00,8'h07,8'h80,8'h1F,8'h00,
8'h07,8'h80,8'h0F,8'h80,8'h07,8'h80,8'h07,8'hC0,8'h07,8'h80,8'h03,8'hC0,8'h07,8'h80,8'h01,8'hE0,
8'h07,8'h80,8'h01,8'hF0,8'h07,8'h80,8'h01,8'hF0,8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h00,8'hF8,
8'h07,8'h80,8'h00,8'hF8,8'h07,8'h80,8'h00,8'hF8,8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,
8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,
8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,
8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,8'h07,8'h80,8'h00,8'h7C,
8'h07,8'h80,8'h00,8'h78,8'h07,8'h80,8'h00,8'hF8,8'h07,8'h80,8'h00,8'hF8,8'h07,8'h80,8'h00,8'hF8,
8'h07,8'h80,8'h00,8'hF0,8'h07,8'h80,8'h01,8'hF0,8'h07,8'h80,8'h01,8'hE0,8'h07,8'h80,8'h03,8'hE0,
8'h07,8'h80,8'h03,8'hC0,8'h07,8'h80,8'h07,8'h80,8'h07,8'h80,8'h1F,8'h80,8'h07,8'h80,8'h3E,8'h00,
8'h0F,8'hC0,8'hFC,8'h00,8'h7F,8'hFF,8'hF0,8'h00,8'h7F,8'hFF,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "D"
    char[40]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h07,8'hE0,8'h00,8'h00,8'h07,8'hE0,8'h00,
8'h00,8'h07,8'hE0,8'h00,8'h00,8'h06,8'hE0,8'h00,8'h00,8'h0C,8'hF0,8'h00,8'h00,8'h0C,8'hF0,8'h00,
8'h00,8'h0C,8'hF0,8'h00,8'h00,8'h0C,8'hF0,8'h00,8'h00,8'h18,8'h78,8'h00,8'h00,8'h18,8'h78,8'h00,
8'h00,8'h18,8'h78,8'h00,8'h00,8'h18,8'h78,8'h00,8'h00,8'h30,8'h3C,8'h00,8'h00,8'h30,8'h3C,8'h00,
8'h00,8'h30,8'h3C,8'h00,8'h00,8'h30,8'h3C,8'h00,8'h00,8'h70,8'h1C,8'h00,8'h00,8'h60,8'h1E,8'h00,
8'h00,8'h60,8'h1E,8'h00,8'h00,8'h60,8'h1E,8'h00,8'h00,8'hE0,8'h0E,8'h00,8'h00,8'hC0,8'h0F,8'h00,
8'h00,8'hC0,8'h0F,8'h00,8'h00,8'hFF,8'hFF,8'h00,8'h01,8'hFF,8'hFF,8'h00,8'h01,8'h80,8'h0F,8'h80,
8'h01,8'h80,8'h07,8'h80,8'h01,8'h80,8'h07,8'h80,8'h03,8'h80,8'h07,8'h80,8'h03,8'h00,8'h07,8'hC0,
8'h03,8'h00,8'h03,8'hC0,8'h03,8'h00,8'h03,8'hC0,8'h07,8'h00,8'h03,8'hC0,8'h06,8'h00,8'h03,8'hE0,
8'h06,8'h00,8'h01,8'hE0,8'h06,8'h00,8'h01,8'hE0,8'h0E,8'h00,8'h01,8'hE0,8'h0E,8'h00,8'h01,8'hF0,
8'h1F,8'h00,8'h01,8'hF8,8'h7F,8'hC0,8'h0F,8'hFE,8'h7F,8'hC0,8'h0F,8'hFE,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "A" 
    char[41]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h0F,8'hFF,8'hFF,8'hF0,8'h0F,8'hFF,8'hFF,8'hF0,8'h0F,8'h03,8'hC0,8'hF8,8'h1E,8'h03,8'hC0,8'h38,
8'h1C,8'h03,8'hC0,8'h38,8'h18,8'h03,8'hC0,8'h18,8'h18,8'h03,8'hC0,8'h18,8'h10,8'h03,8'hC0,8'h0C,
8'h30,8'h03,8'hC0,8'h0C,8'h30,8'h03,8'hC0,8'h04,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,8'h00,8'h03,8'hC0,8'h00,
8'h00,8'h03,8'hE0,8'h00,8'h00,8'h3F,8'hFC,8'h00,8'h00,8'h3F,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "T" 
    char[42]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'hE0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h07,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hF0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h07,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hF0,8'h00,8'h00,8'h00,
8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,
8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h0F,8'hF8,8'h1F,8'hFC,8'h00,8'h00,8'h00,
8'h00,8'h0C,8'h00,8'h3F,8'hFF,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hC0,8'h00,8'h00,
8'h00,8'h00,8'h01,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h00,8'h00,8'h07,8'hFF,8'hF7,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'hE7,8'hF3,8'hFF,8'h00,8'h00,8'h00,8'h00,8'h7F,8'hC7,8'hF0,8'hFF,8'hE0,8'h00,
8'h00,8'h01,8'hFF,8'h87,8'hF0,8'h7F,8'hF8,8'h00,8'h00,8'h0F,8'hFE,8'h03,8'hE0,8'h3F,8'hFF,8'h00,
8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,
8'h3F,8'hFF,8'h9F,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h1F,8'hFE,8'h1F,8'hC0,8'h00,8'hFE,8'h7F,8'hF8,
8'h1F,8'hF8,8'h1F,8'h80,8'h00,8'h7E,8'h3F,8'hF0,8'h07,8'hC0,8'h0F,8'h80,8'h00,8'h7E,8'h0F,8'hE0,
8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFE,8'h03,8'hC0,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFE,8'h00,8'h00,
8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h00,8'h7C,8'h00,8'h00,
8'h00,8'h00,8'h0F,8'h80,8'h00,8'h7C,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,8'h00,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFC,8'h00,8'h00,
8'h00,8'h00,8'h0F,8'hC0,8'h1F,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h06,8'h00,8'h00,8'h70,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'hE0,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,
8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'hFC,8'h00,8'h00,8'h0F,8'hF0,8'h00,8'h00,8'h0F,8'hFC,8'h00,
8'h00,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "查" 
    char[43]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3C,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h07,8'hFE,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7F,8'hFF,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,
8'h00,8'h3F,8'hFF,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h00,8'h07,8'hFF,8'hFF,8'hE0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'hC0,8'h00,8'h00,8'h00,
8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,
8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h03,8'h80,8'h1F,8'h80,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h1F,8'h80,8'h00,8'h00,8'h00,8'h00,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFE,8'h00,
8'h03,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF8,8'h07,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hF0,
8'h0F,8'hFF,8'hC0,8'h3E,8'h00,8'hFF,8'hFF,8'hF0,8'h0F,8'hF8,8'h00,8'h7C,8'h00,8'h01,8'hFF,8'hE0,
8'h0F,8'h00,8'h01,8'hF8,8'h00,8'h00,8'h1F,8'hC0,8'h00,8'h00,8'h03,8'hFF,8'hFF,8'hFF,8'h07,8'h80,
8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'h80,8'h00,
8'h00,8'h00,8'h7F,8'h80,8'h00,8'h3F,8'h80,8'h00,8'h00,8'h01,8'hFF,8'h00,8'h00,8'h3F,8'h80,8'h00,
8'h00,8'h0F,8'hFF,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'h00,8'h7F,8'hFF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,
8'h7F,8'hFF,8'hDF,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h7F,8'hFE,8'h1F,8'h80,8'h00,8'h3F,8'h00,8'h00,
8'h3F,8'hF8,8'h1F,8'h80,8'h00,8'h3F,8'h00,8'h00,8'h1F,8'h80,8'h1F,8'hFF,8'hFF,8'hFF,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'h80,8'h00,8'h3F,8'h00,8'h00,8'h00,8'h00,8'h1F,8'h80,8'h00,8'h3F,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'hFF,8'hF8,8'h3F,8'h00,8'h00,8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'h00,8'h00,8'h00,8'h00,8'h1F,8'hFF,8'hFF,8'hFF,8'h00,8'h00,
8'h00,8'h00,8'h1F,8'h00,8'h00,8'h1E,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "看" 
    char[44]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h80,
8'h00,8'h0F,8'hFF,8'h80,8'h00,8'h00,8'h1F,8'h80,8'h00,8'h0F,8'hFF,8'h8F,8'hFC,8'h00,8'h1F,8'hC0,
8'h00,8'h0F,8'hFF,8'h8F,8'hFE,8'h00,8'h1F,8'hC0,8'h00,8'h0F,8'hFF,8'h9F,8'hFE,8'h00,8'h1F,8'hC0,
8'h00,8'h0F,8'h8F,8'h9F,8'h3E,8'h00,8'h1F,8'hC0,8'h00,8'h0F,8'h8F,8'h9F,8'h3E,8'h06,8'h1F,8'hC0,
8'h00,8'h0F,8'h8F,8'h9F,8'h3E,8'h0F,8'h1F,8'hC0,8'h00,8'h0F,8'h8F,8'h1F,8'h3E,8'h0F,8'h1F,8'hC0,
8'h00,8'h0F,8'h8F,8'h1F,8'h3E,8'h0F,8'h0F,8'hC0,8'h00,8'h0F,8'h8F,8'h1F,8'h3E,8'h0F,8'h0F,8'hC0,
8'h00,8'h0F,8'h8F,8'h1F,8'h3E,8'h0F,8'h0F,8'hC0,8'h00,8'h0F,8'h8F,8'h1F,8'h3E,8'h0F,8'h0F,8'hC0,
8'h0F,8'h0F,8'h8F,8'h1F,8'h3E,8'h0F,8'h0F,8'hC0,8'h1F,8'hFF,8'hFF,8'hFF,8'hFF,8'hCF,8'h0F,8'hC0,
8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hEF,8'h0F,8'hC0,8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hEF,8'h0F,8'hC0,
8'h3F,8'hFF,8'hFF,8'hFF,8'hFF,8'hCF,8'h0F,8'hC0,8'h38,8'h0F,8'h0F,8'h1F,8'h3E,8'h0F,8'h0F,8'hC0,
8'h00,8'h0F,8'h0F,8'h1E,8'h3E,8'h0F,8'h0F,8'hC0,8'h00,8'h0F,8'h0F,8'h1E,8'h3E,8'h0F,8'h0F,8'hC0,
8'h00,8'h0F,8'h0F,8'h1E,8'h3E,8'h0F,8'h0F,8'hC0,8'h00,8'h1F,8'h0F,8'h1E,8'h3E,8'h0F,8'h0F,8'hC0,
8'h00,8'h1F,8'h0F,8'h1E,8'h3E,8'h0F,8'h0F,8'hC0,8'h00,8'h1F,8'h0F,8'h1E,8'h3E,8'h00,8'h1F,8'hC0,
8'h00,8'h3E,8'h0F,8'h1E,8'h3E,8'h00,8'h1F,8'hC0,8'h00,8'h3E,8'h0F,8'h3C,8'h3E,8'h00,8'h1F,8'hC0,
8'h00,8'h7E,8'h0F,8'h3C,8'h3E,8'h00,8'h1F,8'hC0,8'h00,8'h7C,8'h0F,8'h3C,8'h3E,8'h00,8'h1F,8'hC0,
8'h00,8'hFC,8'h0F,8'h78,8'h3E,8'h00,8'h1F,8'hC0,8'h03,8'hF8,8'h0E,8'h78,8'h3E,8'h00,8'h1F,8'hC0,
8'h0F,8'hF8,8'h06,8'hF0,8'h3E,8'h00,8'h3F,8'h80,8'h3F,8'hF0,8'h01,8'hF0,8'h7E,8'h00,8'h7F,8'h80,
8'h3F,8'hE0,8'h07,8'hE0,8'h7E,8'hFF,8'hFF,8'h80,8'h3F,8'h80,8'h0F,8'hC0,8'h3E,8'h7F,8'hFF,8'h80,
8'h0C,8'h00,8'h0F,8'h00,8'h3C,8'h3F,8'hFF,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3C,8'h0F,8'hFE,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "删" 
    char[45]  <= {8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h3C,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7E,8'h00,8'h00,8'h00,
8'h07,8'h00,8'h04,8'h00,8'h7F,8'h00,8'h00,8'h00,8'h0F,8'hFF,8'hFF,8'h00,8'hFE,8'h00,8'h00,8'h00,
8'h3F,8'hFF,8'hFF,8'h01,8'hFF,8'h00,8'h00,8'h00,8'h3F,8'hFF,8'hFF,8'h03,8'hFF,8'hC0,8'h00,8'h00,
8'h3F,8'hFC,8'h7F,8'h07,8'hFF,8'hF8,8'h00,8'h00,8'h11,8'hF0,8'h3E,8'h0F,8'hFF,8'hFE,8'h00,8'h00,
8'h01,8'hF0,8'h3E,8'h0F,8'hE3,8'hFF,8'hE0,8'h00,8'h01,8'hF0,8'h3C,8'h1F,8'h80,8'hFF,8'hFC,8'h00,
8'h01,8'hF0,8'h38,8'h7F,8'h00,8'h7F,8'hFF,8'hC0,8'h01,8'hF0,8'h78,8'hFC,8'h00,8'h1F,8'hFF,8'hFE,
8'h01,8'hF1,8'hF1,8'hF8,8'h00,8'h07,8'hFF,8'hFC,8'h01,8'hFF,8'hF7,8'hE7,8'hF0,8'h03,8'hFF,8'hF8,
8'h01,8'hFF,8'hFF,8'h8F,8'hFF,8'hF8,8'hFF,8'hF8,8'h01,8'hFF,8'hFE,8'h1F,8'hFF,8'hF8,8'h7F,8'hF0,
8'h01,8'hF8,8'h3C,8'h1F,8'hFF,8'h00,8'h1F,8'hE0,8'h01,8'hF8,8'h3C,8'h00,8'h3E,8'h00,8'h07,8'hC0,
8'h01,8'hF8,8'h1C,8'h00,8'h3E,8'h00,8'h00,8'h00,8'h01,8'hF8,8'h1E,8'h3F,8'hFF,8'hFF,8'h00,8'h00,
8'h01,8'hF8,8'h3E,8'h7F,8'hFF,8'hFF,8'h80,8'h00,8'h01,8'hF8,8'h3E,8'hFF,8'hFF,8'hFF,8'hC0,8'h00,
8'h01,8'hF8,8'h7C,8'hFF,8'hFF,8'hFF,8'h80,8'h00,8'h01,8'hF9,8'hFC,8'hF0,8'h3E,8'h00,8'h00,8'h00,
8'h01,8'hFF,8'hF8,8'h00,8'h3E,8'h18,8'h00,8'h00,8'h01,8'hFF,8'hF0,8'h1E,8'h3E,8'h3E,8'h00,8'h00,
8'h01,8'hFF,8'h80,8'h1E,8'h3E,8'h3F,8'h00,8'h00,8'h03,8'hF8,8'h00,8'h3F,8'h3E,8'h3F,8'h80,8'h00,
8'h03,8'hF8,8'h00,8'h7E,8'h3E,8'h3F,8'hC0,8'h00,8'h03,8'hF8,8'h00,8'hFC,8'h3E,8'h1F,8'hE0,8'h00,
8'h03,8'hF8,8'h03,8'hF0,8'h7E,8'h0F,8'hF0,8'h00,8'h03,8'hF0,8'h07,8'hE0,8'h3E,8'h03,8'hF8,8'h00,
8'h03,8'hF0,8'h0F,8'hC0,8'h3E,8'h01,8'hFC,8'h00,8'h03,8'hF0,8'h3F,8'h40,8'h7E,8'h00,8'h7E,8'h00,
8'h03,8'hF0,8'h7C,8'h3F,8'hFF,8'h00,8'h1F,8'h00,8'h03,8'hF0,8'h70,8'h1F,8'hFE,8'h00,8'h03,8'h00,
8'h03,8'hF0,8'h00,8'h0F,8'hFE,8'h00,8'h00,8'h00,8'h03,8'hF0,8'h00,8'h07,8'hFC,8'h00,8'h00,8'h00,
8'h01,8'hE0,8'h00,8'h01,8'hF8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,
8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00} ; // "除"                      

end


// 给不同的界面赋值不同的像素数据
always @(posedge lcd_pclk or negedge sys_rst_n) begin
    if (!sys_rst_n) begin
        pixel_data <= BLACK;
    end else begin
        case (ui_state)
            // 主界面
            2'b00: begin
                // 主界面色块 - 简化优化
                if ((pixel_xpos >= CHAR_POS_X - 1'b1) && (pixel_xpos < CHAR_POS_X + CHAR_WIDTH - 1'b1)
                    && (pixel_ypos >= CHAR_POS_Y) && (pixel_ypos < CHAR_POS_Y + CHAR_HEIGHT)) begin
                    if (char[10][(CHAR_HEIGHT + CHAR_POS_Y - pixel_ypos) * 64 - ((pixel_xpos - (CHAR_POS_X -1'b1)) % 64) - 1'b1])
                        pixel_data <= YELLOW;
                    else
                        pixel_data <= WHITE;
                end
                else if ((pixel_xpos >= CHAR_POS_X + pos_X_remove1 - 1'b1) && (pixel_xpos < CHAR_POS_X + pos_X_remove1 + CHAR_WIDTH - 1'b1)
                    && (pixel_ypos >= CHAR_POS_Y) && (pixel_ypos < CHAR_POS_Y + CHAR_HEIGHT)) begin
                    if (char[11][(CHAR_HEIGHT + CHAR_POS_Y - pixel_ypos) * 64 - ((pixel_xpos - (CHAR_POS_X + pos_X_remove1 -1'b1)) % 64) - 1'b1])
                        pixel_data <= YELLOW;
                    else
                        pixel_data <= WHITE;
                end               
                else if ((pixel_xpos >= CHAR_POS_X + pos_X_remove1*2 - 1'b1) && (pixel_xpos < CHAR_POS_X + pos_X_remove1*2 + CHAR_WIDTH - 1'b1)
                    && (pixel_ypos >= CHAR_POS_Y) && (pixel_ypos < CHAR_POS_Y + CHAR_HEIGHT)) begin
                    if (char[12][(CHAR_HEIGHT + CHAR_POS_Y - pixel_ypos) * 64 - ((pixel_xpos - (CHAR_POS_X + pos_X_remove1*2 -1'b1)) % 64) - 1'b1])
                        pixel_data <= YELLOW;
                    else
                        pixel_data <= WHITE;
                end 
                else if ((pixel_xpos >= CHAR_POS_X + pos_X_remove1*3 - 1'b1) && (pixel_xpos < CHAR_POS_X + pos_X_remove1*3 + CHAR_WIDTH - 1'b1)
                    && (pixel_ypos >= CHAR_POS_Y) && (pixel_ypos < CHAR_POS_Y + CHAR_HEIGHT)) begin
                    if (char[13][(CHAR_HEIGHT + CHAR_POS_Y - pixel_ypos) * 64 - ((pixel_xpos - (CHAR_POS_X + pos_X_remove1*3 -1'b1)) % 64) - 1'b1])
                        pixel_data <= YELLOW;
                    else
                        pixel_data <= WHITE;
                end 
                
                // 心率区域
                else if (pixel_xpos >= xinlv_X_START && pixel_xpos <= xinlv_X_END &&
                    pixel_ypos >= xinlv_Y_START && pixel_ypos <= xinlv_Y_END) begin
                    // 心 (中文64×64)
                    if ((pixel_xpos >= XINLV_TEXT_X - 1'b1) && (pixel_xpos < XINLV_TEXT_X + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= XINLV_TEXT_Y) && (pixel_ypos < XINLV_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[10][(CHINESE_HEIGHT + XINLV_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (XINLV_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(xinlv_bcd_1 > 4'd1 || xinlv_bcd_2 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // 率 (中文64×64)
                    else if ((pixel_xpos >= XINLV_TEXT_X + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < XINLV_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= XINLV_TEXT_Y) && (pixel_ypos < XINLV_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[23][(CHINESE_HEIGHT + XINLV_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (XINLV_TEXT_X + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(xinlv_bcd_1 > 4'd1 || xinlv_bcd_2 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    //心率数据
                    else if ((pixel_xpos >= XINLV_TEXT_X + CHINESE_WIDTH*2+ CHAR_SPACING*2 - 1'b1) && (pixel_xpos < XINLV_TEXT_X +LETTER_WIDTH + CHINESE_WIDTH*2 + CHAR_SPACING*2 - 1'b1)
                        && (pixel_ypos >= XINLV_TEXT_Y) && (pixel_ypos < XINLV_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[xinlv_bcd_1][(CHINESE_HEIGHT + XINLV_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (XINLV_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(xinlv_bcd_1 > 4'd1 || xinlv_bcd_2 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                    else if ((pixel_xpos >= XINLV_TEXT_X + LETTER_WIDTH + CHINESE_WIDTH*2 + CHAR_SPACING*3 - 1'b1) && (pixel_xpos < XINLV_TEXT_X + LETTER_WIDTH*2 + CHINESE_WIDTH*2 + CHAR_SPACING*3 - 1'b1)
                        && (pixel_ypos >= XINLV_TEXT_Y) && (pixel_ypos < XINLV_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[xinlv_bcd_2][(CHINESE_HEIGHT + XINLV_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (XINLV_TEXT_X + LETTER_WIDTH + CHAR_SPACING + CHINESE_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(xinlv_bcd_1 > 4'd1 || xinlv_bcd_2 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                    else if ((pixel_xpos >= XINLV_TEXT_X + LETTER_WIDTH*2 + CHINESE_WIDTH*2 +CHAR_SPACING*4 - 1'b1) && (pixel_xpos < XINLV_TEXT_X + LETTER_WIDTH*3 + CHINESE_WIDTH*2 + CHAR_SPACING*4 - 1'b1)
                        && (pixel_ypos >= XINLV_TEXT_Y) && (pixel_ypos < XINLV_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[xinlv_bcd_3][(CHINESE_HEIGHT + XINLV_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (XINLV_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 + CHINESE_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(xinlv_bcd_1 > 4'd1 || xinlv_bcd_2 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                    else begin
                        if(xinlv_bcd_1 > 4'd1 || xinlv_bcd_2 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                end 
                
                // RR间期区域
                else if (pixel_xpos >= RR_X_START && pixel_xpos <= RR_X_END &&
                    pixel_ypos >= RR_Y_START && pixel_ypos <= RR_Y_END) begin
                    // R (英文32×64)
                    if ((pixel_xpos >= RR_TEXT_X - 1'b1) && (pixel_xpos < RR_TEXT_X + LETTER_WIDTH - 1'b1)
                        && (pixel_ypos >= RR_TEXT_Y) && (pixel_ypos < RR_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[24][(LETTER_HEIGHT + RR_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (RR_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(rr_bcd_1 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // R (英文32×64)
                    else if ((pixel_xpos >= RR_TEXT_X + LETTER_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < RR_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= RR_TEXT_Y) && (pixel_ypos < RR_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[24][(LETTER_HEIGHT + RR_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (RR_TEXT_X + LETTER_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(rr_bcd_1 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // 间 (中文64×64)
                    else if ((pixel_xpos >= RR_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 - 1'b1) && (pixel_xpos < RR_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= RR_TEXT_Y) && (pixel_ypos < RR_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[25][(CHINESE_HEIGHT + RR_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (RR_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(rr_bcd_1 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // 期 (中文64×64)
                    else if ((pixel_xpos >= RR_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < RR_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= RR_TEXT_Y) && (pixel_ypos < RR_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[26][(CHINESE_HEIGHT + RR_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (RR_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(rr_bcd_1 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    //RR间期数据
                    else if ((pixel_xpos >= RR_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 + CHINESE_WIDTH*2 + CHAR_SPACING*2 - 1'b1) && (pixel_xpos < RR_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*2 + CHINESE_WIDTH*2 + CHAR_SPACING*2 - 1'b1)
                        && (pixel_ypos >= RR_TEXT_Y) && (pixel_ypos < RR_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[rr_bcd_1][(CHINESE_HEIGHT + RR_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (RR_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 + CHINESE_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(rr_bcd_1 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                    else if ((pixel_xpos >= RR_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*2 + CHINESE_WIDTH*2 + CHAR_SPACING*3 - 1'b1) && (pixel_xpos < RR_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*2 + CHINESE_WIDTH*2 + CHAR_SPACING*3 - 1'b1)
                        && (pixel_ypos >= RR_TEXT_Y) && (pixel_ypos < RR_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[rr_bcd_2][(CHINESE_HEIGHT + RR_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (RR_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 + CHINESE_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(rr_bcd_1 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                    else if ((pixel_xpos >= RR_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*2 + CHINESE_WIDTH*2 + CHAR_SPACING*4 - 1'b1) && (pixel_xpos < RR_TEXT_X + LETTER_WIDTH*5 + CHAR_SPACING*2 + CHINESE_WIDTH*2 + CHAR_SPACING*4 - 1'b1)
                        && (pixel_ypos >= RR_TEXT_Y) && (pixel_ypos < RR_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[rr_bcd_3][(CHINESE_HEIGHT + RR_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (RR_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 + CHINESE_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(rr_bcd_1 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end

                    else begin
                        if(rr_bcd_1 < 4'd6)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                end 
                
                // HRV区域
                else if (pixel_xpos >= HRV_X_START && pixel_xpos <= HRV_X_END &&
                    pixel_ypos >= HRV_Y_START && pixel_ypos <= HRV_Y_END) begin
                    // H (英文32×64)
                    if ((pixel_xpos >= HRV_TEXT_X - 1'b1) && (pixel_xpos < HRV_TEXT_X + LETTER_WIDTH - 1'b1)
                        && (pixel_ypos >= HRV_TEXT_Y) && (pixel_ypos < HRV_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[27][(LETTER_HEIGHT + HRV_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (HRV_TEXT_X -1'b1)) % 64) - 1'b1])    //设置修改了一下
                            pixel_data <= BLACK;
                        else if(hrv_bcd_2 > 4'd8 || hrv_bcd_2 <4'd2)begin
                            pixel_data <= RED;
                        end
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // R (英文32×64)
                    else if ((pixel_xpos >= HRV_TEXT_X + LETTER_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < HRV_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= HRV_TEXT_Y) && (pixel_ypos < HRV_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[24][(LETTER_HEIGHT + HRV_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (HRV_TEXT_X + LETTER_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(hrv_bcd_2 > 4'd8 || hrv_bcd_2 <4'd2)begin
                            pixel_data <= RED;
                        end
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // V (英文32×64)
                    else if ((pixel_xpos >= HRV_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 - 1'b1) && (pixel_xpos < HRV_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*2 - 1'b1)
                        && (pixel_ypos >= HRV_TEXT_Y) && (pixel_ypos < HRV_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[28][(LETTER_HEIGHT + HRV_TEXT_Y - pixel_ypos) *32 - ((pixel_xpos - (HRV_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(hrv_bcd_2 > 4'd8 || hrv_bcd_2 <4'd2)begin
                            pixel_data <= RED;
                        end
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    //HRV数据
                    else if ((pixel_xpos >= HRV_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 - 1'b1) && (pixel_xpos < HRV_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*3 - 1'b1)
                        && (pixel_ypos >= HRV_TEXT_Y) && (pixel_ypos < HRV_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[hrv_bcd_1][(CHINESE_HEIGHT + HRV_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (HRV_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(hrv_bcd_2 > 4'd8 || hrv_bcd_2 <4'd2)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                    else if ((pixel_xpos >= HRV_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 - 1'b1) && (pixel_xpos < HRV_TEXT_X + LETTER_WIDTH*5 + CHAR_SPACING*4 - 1'b1)
                        && (pixel_ypos >= HRV_TEXT_Y) && (pixel_ypos < HRV_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[hrv_bcd_2][(CHINESE_HEIGHT + HRV_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (HRV_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(hrv_bcd_2 > 4'd8 || hrv_bcd_2 <4'd2)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                    else if ((pixel_xpos >= HRV_TEXT_X + LETTER_WIDTH*5 + CHAR_SPACING*5 - 1'b1) && (pixel_xpos < HRV_TEXT_X + LETTER_WIDTH*6 + CHAR_SPACING*5 - 1'b1)
                        && (pixel_ypos >= HRV_TEXT_Y) && (pixel_ypos < HRV_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[hrv_bcd_3][(CHINESE_HEIGHT + HRV_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (HRV_TEXT_X + LETTER_WIDTH*5 + CHAR_SPACING*5 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else if(hrv_bcd_2 > 4'd8 || hrv_bcd_2 <4'd2)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                    else begin
                        if(hrv_bcd_2 > 4'd8 || hrv_bcd_2 <4'd2)begin
                            pixel_data <= RED;
                        end
                        else begin
                            pixel_data <= LIGHT_GREEN;
                        end
                    end
                end
                    
                // 状态区域
                else if (pixel_xpos >= Level_X_START && pixel_xpos <= Level_X_END &&
                    pixel_ypos >= Level_Y_START && pixel_ypos <= Level_Y_END) begin
                    // 状 (中文64×64)
                    if ((pixel_xpos >= LEVEL_TEXT_X - 1'b1) && (pixel_xpos < LEVEL_TEXT_X + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= LEVEL_TEXT_Y) && (pixel_ypos < LEVEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[29][(CHINESE_HEIGHT + LEVEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (LEVEL_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // 态 (中文64×64)
                    else if ((pixel_xpos >= LEVEL_TEXT_X + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < LEVEL_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= LEVEL_TEXT_Y) && (pixel_ypos < LEVEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[30][(CHINESE_HEIGHT + LEVEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (LEVEL_TEXT_X + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    //状态文字
                    else if ((pixel_xpos >= LEVEL_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING*2 - 1'b1) && (pixel_xpos < LEVEL_TEXT_X + CHINESE_WIDTH*3 + CHAR_SPACING*2 - 1'b1)
                        && (pixel_ypos >= LEVEL_TEXT_Y) && (pixel_ypos < LEVEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[level_state[0]][(CHINESE_HEIGHT + LEVEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (LEVEL_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    else if ((pixel_xpos >= LEVEL_TEXT_X + CHINESE_WIDTH*3 + CHAR_SPACING*3 - 1'b1) && (pixel_xpos < LEVEL_TEXT_X + CHINESE_WIDTH*4 + CHAR_SPACING*3 - 1'b1)
                        && (pixel_ypos >= LEVEL_TEXT_Y) && (pixel_ypos < LEVEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[level_state[1]][(CHINESE_HEIGHT + LEVEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (LEVEL_TEXT_X + CHINESE_WIDTH*3 + CHAR_SPACING*3 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end

                    /*
                    else if ((pixel_xpos >= LEVEL_TEXT_X + CHINESE_WIDTH*4 + CHAR_SPACING*4 - 1'b1) && (pixel_xpos < LEVEL_TEXT_X + CHINESE_WIDTH*5 + CHAR_SPACING*4 - 1'b1)
                        && (pixel_ypos >= LEVEL_TEXT_Y) && (pixel_ypos < LEVEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[level_state[3]][(CHINESE_HEIGHT + LEVEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (LEVEL_TEXT_X + CHINESE_WIDTH*4 + CHAR_SPACING*4 -1'b1)) % 64) - 1'b1] && arrhythmia_level != 2'd0)
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    else if ((pixel_xpos >= LEVEL_TEXT_X + CHINESE_WIDTH*5 + CHAR_SPACING*5 - 1'b1) && (pixel_xpos < LEVEL_TEXT_X + CHINESE_WIDTH*6 + CHAR_SPACING*5 - 1'b1)
                        && (pixel_ypos >= LEVEL_TEXT_Y) && (pixel_ypos < LEVEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[level_state[4]][(CHINESE_HEIGHT + LEVEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (LEVEL_TEXT_X + CHINESE_WIDTH*5 + CHAR_SPACING*5 -1'b1)) % 64) - 1'b1] && arrhythmia_level != 2'd0)
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN  
                    end
                    */
                    else begin
                        pixel_data <= LIGHT_GREEN;
                    end
                end 

                // 心电图按钮
                else if (pixel_xpos >= xdt_X_START && pixel_xpos <= xdt_X_END &&
                    pixel_ypos >= xdt_Y_START && pixel_ypos <= xdt_Y_END) begin
                    // 按钮边框
                    if (pixel_xpos == xdt_X_START || pixel_xpos == xdt_X_END ||
                        pixel_ypos == xdt_Y_START || pixel_ypos == xdt_Y_END) begin
                        pixel_data <= BLACK;
                    end 
                    // 心 (中文64×64)
                    else if ((pixel_xpos >= XDT_TEXT_X - 1'b1) && (pixel_xpos < XDT_TEXT_X + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= XDT_TEXT_Y) && (pixel_ypos < XDT_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[10][(CHINESE_HEIGHT + XDT_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (XDT_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 电 (中文64×64)
                    else if ((pixel_xpos >= XDT_TEXT_X + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < XDT_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= XDT_TEXT_Y) && (pixel_ypos < XDT_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[14][(CHINESE_HEIGHT + XDT_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (XDT_TEXT_X + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 波 (中文64×64)
                    else if ((pixel_xpos >= XDT_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING*2 - 1'b1) && (pixel_xpos < XDT_TEXT_X + CHINESE_WIDTH*3 + CHAR_SPACING*2 - 1'b1)
                        && (pixel_ypos >= XDT_TEXT_Y) && (pixel_ypos < XDT_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[15][(CHINESE_HEIGHT + XDT_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (XDT_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    //形
                    else if ((pixel_xpos >= XDT_TEXT_X + CHINESE_WIDTH*3 + CHAR_SPACING*3 - 1'b1) && (pixel_xpos < XDT_TEXT_X + CHINESE_WIDTH*4 + CHAR_SPACING*3 - 1'b1)
                        && (pixel_ypos >= XDT_TEXT_Y) && (pixel_ypos < XDT_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[16][(CHINESE_HEIGHT + XDT_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (XDT_TEXT_X + CHINESE_WIDTH*3 + CHAR_SPACING*3 -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 按钮内部
                    else begin
                        pixel_data <= LIGHT_BLUE;
                    end
                end 
                
                // 心率回看按钮
                else if (pixel_xpos >= save_X_START && pixel_xpos <= save_X_END &&
                         pixel_ypos >= save_Y_START && pixel_ypos <= save_Y_END) begin
                    // 按钮边框
                    if (pixel_xpos == save_X_START || pixel_xpos == save_X_END ||
                        pixel_ypos == save_Y_START || pixel_ypos == save_Y_END) begin
                        pixel_data <= BLACK;
                    end 
                    // 记 (中文64×64)
                    else if ((pixel_xpos >= SAVE_TEXT_X - 1'b1) && (pixel_xpos < SAVE_TEXT_X + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= SAVE_TEXT_Y) && (pixel_ypos < SAVE_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[17][(CHINESE_HEIGHT + SAVE_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (SAVE_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 录 (中文64×64)
                    else if ((pixel_xpos >= SAVE_TEXT_X + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < SAVE_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= SAVE_TEXT_Y) && (pixel_ypos < SAVE_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[18][(CHINESE_HEIGHT + SAVE_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (SAVE_TEXT_X + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 按钮内部
                    else begin
                        pixel_data <= LIGHT_BLUE;
                    end
                end

                // 搜索按钮
                else if (pixel_xpos >= search_X_START && pixel_xpos <= search_X_END &&
                         pixel_ypos >= search_Y_START && pixel_ypos <= search_Y_END) begin
                    // 按钮边框
                    if (pixel_xpos == search_X_START || pixel_xpos == search_X_END ||
                        pixel_ypos == search_Y_START || pixel_ypos == search_Y_END) begin
                        pixel_data <= BLACK;
                    end 
                    // 检 (中文64×64)
                    else if ((pixel_xpos >= SEARCH_TEXT_X - 1'b1) && (pixel_xpos < SEARCH_TEXT_X + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= SEARCH_TEXT_Y) && (pixel_ypos < SEARCH_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[19][(CHINESE_HEIGHT + SEARCH_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (SEARCH_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 索 (中文64×64)
                    else if ((pixel_xpos >= SEARCH_TEXT_X + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < SEARCH_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= SEARCH_TEXT_Y) && (pixel_ypos < SEARCH_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[20][(CHINESE_HEIGHT + SEARCH_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (SEARCH_TEXT_X + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 按钮内部
                    else begin
                        pixel_data <= LIGHT_BLUE;
                    end
                end

                else begin
                    // 背景
                    pixel_data <= WHITE;
                end
            end
            
            // 心电图显示界面
            2'b01: begin
                // 返回按钮
                if (pixel_xpos >= return_X_START && pixel_xpos <= return_X_END &&
                    pixel_ypos >= return_Y_START && pixel_ypos <= return_Y_END) begin
                    // 按钮边框
                    if (pixel_xpos == return_X_START || pixel_xpos == return_X_END ||
                        pixel_ypos == return_Y_START || pixel_ypos == return_Y_END) begin
                        pixel_data <= BLACK;
                    end 
                    // 返 (中文64×64)
                    else if ((pixel_xpos >= RETURN_TEXT_X - 1'b1) && (pixel_xpos < RETURN_TEXT_X + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= RETURN_TEXT_Y) && (pixel_ypos < RETURN_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[21][(CHINESE_HEIGHT + RETURN_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (RETURN_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= RED;
                    end
                    // 回 (中文64×64)
                    else if ((pixel_xpos >= RETURN_TEXT_X + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < RETURN_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= RETURN_TEXT_Y) && (pixel_ypos < RETURN_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[22][(CHINESE_HEIGHT + RETURN_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (RETURN_TEXT_X + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= RED;
                    end
                    // 按钮内部
                    else begin
                        pixel_data <= RED;
                    end
                end
                else begin
                    // 背景
                    pixel_data <= WHITE;
                end
            end
            
            // 心率回看界面
            2'b10: begin
                // 返回按钮
                if (pixel_xpos >= return_X_START && pixel_xpos <= return_X_END &&
                    pixel_ypos >= return_Y_START && pixel_ypos <= return_Y_END) begin
                    // 按钮边框
                    if (pixel_xpos == return_X_START || pixel_xpos == return_X_END ||
                        pixel_ypos == return_Y_START || pixel_ypos == return_Y_END) begin
                        pixel_data <= BLACK;
                    end 
                    // 返 (中文64×64)
                    else if ((pixel_xpos >= RETURN_TEXT_X - 1'b1) && (pixel_xpos < RETURN_TEXT_X + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= RETURN_TEXT_Y) && (pixel_ypos < RETURN_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[21][(CHINESE_HEIGHT + RETURN_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (RETURN_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= RED;
                    end
                    // 回 (中文64×64)
                    else if ((pixel_xpos >= RETURN_TEXT_X + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < RETURN_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= RETURN_TEXT_Y) && (pixel_ypos < RETURN_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[22][(CHINESE_HEIGHT + RETURN_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (RETURN_TEXT_X + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= RED;
                    end
                    // 按钮内部
                    else begin
                        pixel_data <= RED;
                    end
                end

                // 选择按钮
                else if (pixel_xpos >= sel_X_START && pixel_xpos <= sel_X_END &&
                    pixel_ypos >= sel_Y_START && pixel_ypos <= sel_Y_END) begin
                    // 按钮边框
                    if (pixel_xpos == sel_X_START || pixel_xpos == sel_X_END ||
                        pixel_ypos == sel_Y_START || pixel_ypos == sel_Y_END) begin
                        pixel_data <= BLACK;
                    end 
                    // 选 (中文64×64)
                    else if ((pixel_xpos >= SEL_TEXT_X - 1'b1) && (pixel_xpos < SEL_TEXT_X + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= SEL_TEXT_Y) && (pixel_ypos < SEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[42][(CHINESE_HEIGHT + SEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (SEL_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 择 (中文64×64)
                    else if ((pixel_xpos >= SEL_TEXT_X + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < SEL_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= SEL_TEXT_Y) && (pixel_ypos < SEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[43][(CHINESE_HEIGHT + SEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (SEL_TEXT_X + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 按钮内部
                    else begin
                        pixel_data <= LIGHT_BLUE;
                    end
                end

                // 删除按钮
                else if (pixel_xpos >= del_X_START && pixel_xpos <= del_X_END &&
                    pixel_ypos >= del_Y_START && pixel_ypos <= del_Y_END) begin
                    // 按钮边框
                    if (pixel_xpos == del_X_START || pixel_xpos == del_X_END ||
                        pixel_ypos == del_Y_START || pixel_ypos == del_Y_END) begin
                        pixel_data <= BLACK;
                    end 
                    // 删 (中文64×64)
                    else if ((pixel_xpos >= DEL_TEXT_X - 1'b1) && (pixel_xpos < DEL_TEXT_X + CHINESE_WIDTH - 1'b1)
                        && (pixel_ypos >= DEL_TEXT_Y) && (pixel_ypos < DEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[44][(CHINESE_HEIGHT + DEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (DEL_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 除 (中文64×64)
                    else if ((pixel_xpos >= DEL_TEXT_X + CHINESE_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < DEL_TEXT_X + CHINESE_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= DEL_TEXT_Y) && (pixel_ypos < DEL_TEXT_Y + CHINESE_HEIGHT)) begin
                        if (char[45][(CHINESE_HEIGHT + DEL_TEXT_Y - pixel_ypos) * 64 - ((pixel_xpos - (DEL_TEXT_X + CHINESE_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= GRAY;
                        else
                            pixel_data <= LIGHT_BLUE;
                    end
                    // 按钮内部
                    else begin
                        pixel_data <= LIGHT_BLUE;
                    end
                end
                
                // 数据选择色块 - DATA1
                else if (pixel_xpos >= data1_X_START && pixel_xpos <= data1_X_END &&
                    pixel_ypos >= data1_Y_START && pixel_ypos <= data1_Y_END && data_state > 3'd0) begin
                    // D (英文32×64)
                    if ((pixel_xpos >= DATA1_TEXT_X - 1'b1) && (pixel_xpos < DATA1_TEXT_X + LETTER_WIDTH - 1'b1)
                        && (pixel_ypos >= DATA1_TEXT_Y) && (pixel_ypos < DATA1_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[39][(LETTER_HEIGHT + DATA1_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA1_TEXT_X -1'b1)) % 32) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // A (英文32×64)
                    else if ((pixel_xpos >= DATA1_TEXT_X + LETTER_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < DATA1_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= DATA1_TEXT_Y) && (pixel_ypos < DATA1_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[40][(LETTER_HEIGHT + DATA1_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA1_TEXT_X + LETTER_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // T (英文32×64)
                    else if ((pixel_xpos >= DATA1_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 - 1'b1) && (pixel_xpos < DATA1_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*2 - 1'b1)
                        && (pixel_ypos >= DATA1_TEXT_Y) && (pixel_ypos < DATA1_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[41][(LETTER_HEIGHT + DATA1_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA1_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // A (英文32×64)
                    else if ((pixel_xpos >= DATA1_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 - 1'b1) && (pixel_xpos < DATA1_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*3 - 1'b1)
                        && (pixel_ypos >= DATA1_TEXT_Y) && (pixel_ypos < DATA1_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[40][(LETTER_HEIGHT + DATA1_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA1_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // 1 (英文32×64)
                    else if ((pixel_xpos >= DATA1_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 - 1'b1) && (pixel_xpos < DATA1_TEXT_X + LETTER_WIDTH*5 + CHAR_SPACING*4 - 1'b1)
                        && (pixel_ypos >= DATA1_TEXT_Y) && (pixel_ypos < DATA1_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[1][(LETTER_HEIGHT + DATA1_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA1_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    else begin
                        pixel_data <= LIGHT_GREEN;
                    end
                end 
                
                // 数据选择色块 - DATA2
                else if (pixel_xpos >= data2_X_START && pixel_xpos <= data2_X_END &&
                    pixel_ypos >= data2_Y_START && pixel_ypos <= data2_Y_END && data_state > 3'd1) begin
                    // D (英文32×64)
                    if ((pixel_xpos >= DATA2_TEXT_X - 1'b1) && (pixel_xpos < DATA2_TEXT_X + LETTER_WIDTH - 1'b1)
                        && (pixel_ypos >= DATA2_TEXT_Y) && (pixel_ypos < DATA2_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[39][(LETTER_HEIGHT + DATA2_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA2_TEXT_X -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // A (英文32×64)
                    else if ((pixel_xpos >= DATA2_TEXT_X + LETTER_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < DATA2_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= DATA2_TEXT_Y) && (pixel_ypos < DATA2_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[40][(LETTER_HEIGHT + DATA2_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA2_TEXT_X + LETTER_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // T (英文32×64)
                    else if ((pixel_xpos >= DATA2_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 - 1'b1) && (pixel_xpos < DATA2_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*2 - 1'b1)
                        && (pixel_ypos >= DATA2_TEXT_Y) && (pixel_ypos < DATA2_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[41][(LETTER_HEIGHT + DATA2_TEXT_Y - pixel_ypos) * 32- ((pixel_xpos - (DATA2_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // A (英文32×64)
                    else if ((pixel_xpos >= DATA2_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 - 1'b1) && (pixel_xpos < DATA2_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*3 - 1'b1)
                        && (pixel_ypos >= DATA2_TEXT_Y) && (pixel_ypos < DATA2_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[40][(LETTER_HEIGHT + DATA2_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA2_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // 2 (英文32×64)
                    else if ((pixel_xpos >= DATA2_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 - 1'b1) && (pixel_xpos < DATA2_TEXT_X + LETTER_WIDTH*5 + CHAR_SPACING*4 - 1'b1)
                        && (pixel_ypos >= DATA2_TEXT_Y) && (pixel_ypos < DATA2_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[2][(LETTER_HEIGHT + DATA2_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA2_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    else begin
                        pixel_data <= LIGHT_GREEN;
                    end
                end 
                
                // 数据选择色块 - DATA3
                else if (pixel_xpos >= data3_X_START && pixel_xpos <= data3_X_END &&
                    pixel_ypos >= data3_Y_START && pixel_ypos <= data3_Y_END && data_state > 3'd2) begin
                    // D (英文32×64)
                    if ((pixel_xpos >= DATA3_TEXT_X - 1'b1) && (pixel_xpos < DATA3_TEXT_X + LETTER_WIDTH - 1'b1)
                        && (pixel_ypos >= DATA3_TEXT_Y) && (pixel_ypos < DATA3_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[39][(LETTER_HEIGHT + DATA3_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA3_TEXT_X -1'b1)) % 32) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // A (英文32×64)
                    else if ((pixel_xpos >= DATA3_TEXT_X + LETTER_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < DATA3_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= DATA3_TEXT_Y) && (pixel_ypos < DATA3_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[40][(LETTER_HEIGHT + DATA3_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA3_TEXT_X + LETTER_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // T (英文32×64)
                    else if ((pixel_xpos >= DATA3_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 - 1'b1) && (pixel_xpos < DATA3_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*2 - 1'b1)
                        && (pixel_ypos >= DATA3_TEXT_Y) && (pixel_ypos < DATA3_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[41][(LETTER_HEIGHT + DATA3_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA3_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // A (英文32×64)
                    else if ((pixel_xpos >= DATA3_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 - 1'b1) && (pixel_xpos < DATA3_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*3 - 1'b1)
                        && (pixel_ypos >= DATA3_TEXT_Y) && (pixel_ypos < DATA3_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[40][(LETTER_HEIGHT + DATA3_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA3_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // 3 (英文32×64)
                    else if ((pixel_xpos >= DATA3_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 - 1'b1) && (pixel_xpos < DATA3_TEXT_X + LETTER_WIDTH*5 + CHAR_SPACING*4 - 1'b1)
                        && (pixel_ypos >= DATA3_TEXT_Y) && (pixel_ypos < DATA3_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[3][(LETTER_HEIGHT + DATA3_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA3_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    else begin
                        pixel_data <= LIGHT_GREEN;
                    end
                end 
                
                // 数据选择色块 - DATA4
                else if (pixel_xpos >= data4_X_START && pixel_xpos <= data4_X_END &&
                    pixel_ypos >= data4_Y_START && pixel_ypos <= data4_Y_END && data_state > 3'd3) begin
                    // D (英文32×64)
                    if ((pixel_xpos >= DATA4_TEXT_X - 1'b1) && (pixel_xpos < DATA4_TEXT_X + LETTER_WIDTH - 1'b1)
                        && (pixel_ypos >= DATA4_TEXT_Y) && (pixel_ypos < DATA4_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[39][(LETTER_HEIGHT + DATA4_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA4_TEXT_X -1'b1)) % 32) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // A (英文32×64)
                    else if ((pixel_xpos >= DATA4_TEXT_X + LETTER_WIDTH + CHAR_SPACING - 1'b1) && (pixel_xpos < DATA4_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING - 1'b1)
                        && (pixel_ypos >= DATA4_TEXT_Y) && (pixel_ypos < DATA4_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[40][(LETTER_HEIGHT + DATA4_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA4_TEXT_X + LETTER_WIDTH + CHAR_SPACING -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // T (英文32×64)
                    else if ((pixel_xpos >= DATA4_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 - 1'b1) && (pixel_xpos < DATA4_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*2 - 1'b1)
                        && (pixel_ypos >= DATA4_TEXT_Y) && (pixel_ypos < DATA4_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[41][(LETTER_HEIGHT + DATA4_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA4_TEXT_X + LETTER_WIDTH*2 + CHAR_SPACING*2 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // A (英文32×64)
                    else if ((pixel_xpos >= DATA4_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 - 1'b1) && (pixel_xpos < DATA4_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*3 - 1'b1)
                        && (pixel_ypos >= DATA4_TEXT_Y) && (pixel_ypos < DATA4_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[40][(LETTER_HEIGHT + DATA4_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA4_TEXT_X + LETTER_WIDTH*3 + CHAR_SPACING*3 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    // 4 (英文32×64)
                    else if ((pixel_xpos >= DATA4_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 - 1'b1) && (pixel_xpos < DATA4_TEXT_X + LETTER_WIDTH*5 + CHAR_SPACING*4 - 1'b1)
                        && (pixel_ypos >= DATA4_TEXT_Y) && (pixel_ypos < DATA4_TEXT_Y + LETTER_HEIGHT)) begin
                        if (char[4][(LETTER_HEIGHT + DATA4_TEXT_Y - pixel_ypos) * 32 - ((pixel_xpos - (DATA4_TEXT_X + LETTER_WIDTH*4 + CHAR_SPACING*4 -1'b1)) % 64) - 1'b1])
                            pixel_data <= BLACK;
                        else
                            pixel_data <= LIGHT_GREEN;
                    end
                    else begin
                        pixel_data <= LIGHT_GREEN;
                    end
                end 

                else begin
                    // 背景
                    pixel_data <= WHITE;
                end
            end
            
            default: pixel_data <= WHITE;
        endcase
    end
end

endmodule